netcdf file\:/home/walter/TechX/ceres/datasets/GLASS {
  dimensions:
    time = 2693;
  variables:
    int base_time;
      base_time:long_name = "sounding launch time";
      base_time:units = "seconds since 1970-01-01 00:00:00 UTC";
      base_time:string = "Fri Jun 30 00:49:09 2000";

    float time_offset(time);
      time_offset:long_name = "seconds since base_time";
      time_offset:units = "seconds";
      time_offset:missing_value = -999.0f;
      time_offset:_FillValue = -999.0f;

    double time(time);
      time:long_name = "time";
      time:units = "seconds since 1970-01-01 00:00:00 UTC";
      time:missing_value = -999.0f;
      time:_FillValue = -999.0;

    float pres(time);
      pres:long_name = "pres";
      pres:units = "mb";
      pres:missing_value = -999.0f;
      pres:_FillValue = -999.0f;

    float tdry(time);
      tdry:long_name = "tdry";
      tdry:units = "deg C";
      tdry:missing_value = -999.0f;
      tdry:_FillValue = -999.0f;

    float dp(time);
      dp:long_name = "dp";
      dp:units = "deg C";
      dp:missing_value = -999.0f;
      dp:_FillValue = -999.0f;

    float rh(time);
      rh:long_name = "rh";
      rh:units = "percent";
      rh:missing_value = -999.0f;
      rh:_FillValue = -999.0f;

    float u_wind(time);
      u_wind:long_name = "u_wind";
      u_wind:units = "m/s";
      u_wind:missing_value = -999.0f;
      u_wind:_FillValue = -999.0f;

    float v_wind(time);
      v_wind:long_name = "v_wind";
      v_wind:units = "m/s";
      v_wind:missing_value = -999.0f;
      v_wind:_FillValue = -999.0f;

    float wspd(time);
      wspd:long_name = "wspd";
      wspd:units = "m/s";
      wspd:missing_value = -999.0f;
      wspd:_FillValue = -999.0f;

    float wdir(time);
      wdir:long_name = "wdir";
      wdir:units = "degree";
      wdir:missing_value = -999.0f;
      wdir:_FillValue = -999.0f;

    float dz(time);
      dz:long_name = "dz";
      dz:units = "m/s";
      dz:missing_value = -999.0f;
      dz:_FillValue = -999.0f;

    float range(time);
      range:long_name = "range";
      range:units = "km";
      range:missing_value = -999.0f;
      range:_FillValue = -999.0f;

    float qp(time);
      qp:long_name = "qp";
      qp:units = "mb";
      qp:missing_value = -999.0f;
      qp:_FillValue = -999.0f;

    float qt(time);
      qt:long_name = "qt";
      qt:units = "deg C";
      qt:missing_value = -999.0f;
      qt:_FillValue = -999.0f;

    float qrh(time);
      qrh:long_name = "qrh";
      qrh:units = "percent";
      qrh:missing_value = -999.0f;
      qrh:_FillValue = -999.0f;

    float qu(time);
      qu:long_name = "qu";
      qu:units = "m/s";
      qu:missing_value = -999.0f;
      qu:_FillValue = -999.0f;

    float qv(time);
      qv:long_name = "qv";
      qv:units = "m/s";
      qv:missing_value = -999.0f;
      qv:_FillValue = -999.0f;

    float qwind(time);
      qwind:long_name = "qwind";
      qwind:units = "m/s";
      qwind:missing_value = -999.0f;
      qwind:_FillValue = -999.0f;

    float mr(time);
      mr:long_name = "mr";
      mr:units = "g/kg";
      mr:missing_value = -999.0f;
      mr:_FillValue = -999.0f;

    float vt(time);
      vt:long_name = "vt";
      vt:units = "deg C";
      vt:missing_value = -999.0f;
      vt:_FillValue = -999.0f;

    float theta(time);
      theta:long_name = "theta";
      theta:units = "deg K";
      theta:missing_value = -999.0f;
      theta:_FillValue = -999.0f;

    float theta_e(time);
      theta_e:long_name = "theta_e";
      theta_e:units = "deg K";
      theta_e:missing_value = -999.0f;
      theta_e:_FillValue = -999.0f;

    float theta_v(time);
      theta_v:long_name = "theta_v";
      theta_v:units = "deg K";
      theta_v:missing_value = -999.0f;
      theta_v:_FillValue = -999.0f;

    float lat(time);
      lat:long_name = "north latitude";
      lat:units = "degrees";
      lat:missing_value = -999.0f;
      lat:_FillValue = -999.0f;
      lat:valid_range = -90.0f, 90.0f;

    float lon(time);
      lon:long_name = "east longitude";
      lon:units = "degrees";
      lon:missing_value = -999.0f;
      lon:_FillValue = -999.0f;
      lon:valid_range = -180.0f, 180.0f;

    float alt(time);
      alt:long_name = "altitude";
      alt:units = "meters";
      alt:missing_value = -999.0f;
      alt:_FillValue = -999.0f;

  // global attributes:
  :bad_value_flag = -999.0f;
  :zebra_platform = "class";
  :history = "ClassNcFile";
  :AvapsEditorVersion = "2.2.2";
  :SoundingDescription = "D200006292355.st1 Version:       STEPS Mobile 1, GLASS 2.01\r  ";
  :ACagency = "AF001";
  :ACtype = "0";
  :AbrHdrOvr = "";
  :BaudRateIndex = "2";
  :CommPortIndex = "0";
  :IcaoIndex = "1";
  :MissionId = "TRAIN";
  :MissionStorm = "WXWXA";
  :OptIcao = "";
  :OptionAutoFile = "1";
  :OptionBSN = "99999";
  :OptionCallSign = "CALL";
  :OptionChuteArea = "676";
  :OptionDoLevels = "1";
  :OptionDoQC = "1";
  :OptionDoWMO = "1";
  :OptionDropSondeMass = "395";
  :OptionPosInterpSpan = "60";
  :OptionTempMsgType = "2";
  :PresBuddySlope = "2";
  :PresOffset = "0";
  :PresOutlier = "10";
  :PresQCDev = "3";
  :PresQCWL = "60";
  :PresSmoothWL = "60";
  :QCSaveDir = "H:\\steps";
  :RHBuddySlope = "20";
  :RHOffset = "0";
  :RHOutlier = "10";
  :RHQCDev = "3";
  :RHQCWL = "60";
  :RHSmoothWL = "60";
  :RawSaveDir = "";
  :SfcAltUnknown = "0";
  :SfcAltitude = "955.1";
  :TdryBuddySlope = "3";
  :TdryDynCor = "1";
  :TdryOffset = "0";
  :TdryOutlier = "10";
  :TdryQCDev = "3";
  :TdryQCWL = "60";
  :TdrySmoothWL = "60";
  :WindBuddySlope = "5";
  :WindDynCor = "1";
  :WindOutlier = "10";
  :WindQCDev = "3";
  :WindQCWL = "10";
  :WindSats = "3";
  :WindSmoothWL = "10";
  :WindVVdelta = "2.5";
  :WmoSaveDir = "C:\\";
  :excludeAbrHdr = "0";
 data:
base_time =962347749
time_offset =
  {-1.0, 0.0, 1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0, 51.0, 52.0, 53.0, 54.0, 55.0, 56.0, 57.0, 58.0, 59.1, 60.1, 61.1, 62.1, 63.1, 64.1, 65.1, 66.1, 67.1, 68.1, 69.1, 70.1, 71.1, 72.1, 73.1, 74.1, 75.1, 76.1, 77.1, 78.1, 79.1, 80.1, 81.1, 82.1, 83.1, 84.1, 85.1, 86.1, 87.1, 88.1, 89.1, 90.1, 91.1, 92.1, 93.1, 94.1, 95.1, 96.1, 97.1, 98.1, 99.1, 100.1, 101.1, 102.1, 103.1, 104.1, 105.1, 106.1, 107.1, 108.1, 109.1, 110.1, 111.1, 112.1, 113.1, 114.1, 115.1, 116.1, 117.1, 118.1, 119.1, 120.1, 121.1, 122.1, 123.1, 124.1, 125.1, 126.1, 127.1, 128.1, 129.1, 130.1, 131.1, 132.1, 133.1, 134.1, 135.1, 136.1, 137.1, 138.1, 139.1, 140.1, 141.1, 142.1, 143.1, 144.1, 145.1, 146.1, 147.1, 148.1, 149.1, 150.1, 151.1, 152.1, 153.1, 154.1, 155.1, 156.1, 157.1, 158.2, 159.2, 160.2, 161.2, 162.2, 163.2, 164.2, 165.2, 166.2, 167.2, 168.2, 169.2, 170.2, 171.2, 172.2, 173.2, 174.2, 175.2, 176.2, 177.2, 178.2, 179.2, 180.2, 181.2, 182.2, 183.2, 184.2, 185.2, 186.2, 187.2, 188.2, 189.2, 190.2, 191.2, 192.2, 193.2, 194.2, 195.2, 196.2, 197.2, 198.2, 199.2, 200.2, 201.2, 202.2, 203.2, 204.2, 205.2, 206.2, 207.2, 208.2, 209.2, 210.2, 211.2, 212.2, 213.2, 214.2, 215.2, 216.2, 217.2, 218.2, 219.2, 220.2, 221.2, 222.2, 223.2, 224.2, 225.2, 226.2, 227.2, 228.2, 229.2, 230.2, 231.2, 232.2, 233.2, 234.2, 235.2, 236.2, 237.2, 238.2, 239.2, 240.2, 241.2, 242.2, 243.2, 244.2, 245.2, 246.2, 247.2, 248.2, 249.2, 250.2, 251.2, 252.2, 253.2, 254.2, 255.2, 256.2, 257.2, 258.2, 259.2, 260.2, 261.2, 262.3, 263.3, 264.3, 265.3, 266.3, 267.3, 268.3, 269.3, 270.3, 271.3, 272.3, 273.3, 274.3, 275.3, 276.3, 277.3, 278.3, 279.3, 280.3, 281.3, 282.3, 283.3, 284.3, 285.3, 286.3, 287.3, 288.3, 289.3, 290.3, 291.3, 292.3, 293.3, 294.3, 295.3, 296.3, 297.3, 298.3, 299.3, 300.3, 301.3, 302.3, 303.3, 304.3, 305.3, 306.3, 307.3, 308.3, 309.3, 310.3, 311.3, 312.3, 313.3, 314.3, 315.3, 316.3, 317.3, 318.3, 319.3, 320.3, 321.3, 322.3, 323.3, 324.3, 325.3, 326.3, 327.3, 328.3, 329.3, 330.3, 331.3, 332.3, 333.3, 334.3, 335.3, 336.3, 337.3, 338.3, 339.3, 340.3, 341.3, 342.3, 343.3, 344.3, 345.3, 346.3, 347.3, 348.3, 349.3, 350.3, 351.3, 352.3, 353.3, 354.3, 355.3, 356.3, 357.3, 358.3, 359.3, 360.3, 361.3, 362.3, 363.3, 364.4, 365.4, 366.4, 367.4, 368.4, 369.4, 370.4, 371.4, 372.4, 373.4, 374.4, 375.4, 376.4, 377.4, 378.4, 379.4, 380.4, 381.4, 382.4, 383.4, 384.4, 385.4, 386.4, 387.4, 388.4, 389.4, 390.4, 391.4, 392.4, 393.4, 394.4, 395.4, 396.4, 397.4, 398.4, 399.4, 400.4, 401.4, 402.4, 403.4, 404.4, 405.4, 406.4, 407.4, 408.4, 409.4, 410.4, 411.4, 412.4, 413.4, 414.4, 415.4, 416.4, 417.4, 418.4, 419.4, 420.4, 421.4, 422.4, 423.4, 424.4, 425.4, 426.4, 427.4, 428.4, 429.4, 430.4, 431.4, 432.4, 433.4, 434.4, 435.4, 436.4, 437.4, 438.4, 439.4, 440.4, 441.4, 442.4, 443.4, 444.4, 445.4, 446.4, 447.4, 448.4, 449.4, 450.4, 451.4, 452.4, 453.4, 454.4, 455.4, 456.5, 457.5, 458.5, 459.5, 460.5, 461.5, 462.5, 463.5, 464.5, 465.5, 466.5, 467.5, 468.5, 469.5, 470.5, 471.5, 472.5, 473.5, 474.5, 475.5, 476.5, 477.5, 478.5, 479.5, 480.5, 481.5, 482.5, 483.5, 484.5, 485.5, 486.5, 487.5, 488.5, 489.5, 490.5, 491.5, 492.5, 493.5, 494.5, 495.5, 496.5, 497.5, 498.5, 499.5, 500.5, 501.5, 502.5, 503.5, 504.5, 505.5, 506.5, 507.5, 508.5, 509.5, 510.5, 511.5, 512.5, 513.5, 514.5, 515.5, 516.5, 517.5, 518.5, 519.5, 520.5, 521.5, 522.5, 523.5, 524.5, 525.5, 526.5, 527.5, 528.5, 529.5, 530.5, 531.5, 532.5, 533.5, 534.5, 535.5, 536.5, 537.5, 538.5, 539.5, 540.5, 541.5, 542.5, 543.5, 544.5, 545.5, 546.5, 547.5, 548.5, 549.5, 550.5, 551.5, 552.5, 553.5, 554.5, 555.5, 556.5, 557.5, 558.5, 559.5, 560.5, 561.5, 562.5, 563.5, 564.5, 565.5, 566.5, 567.5, 568.6, 569.6, 570.6, 571.6, 572.6, 573.6, 574.6, 575.6, 576.6, 577.6, 578.6, 579.6, 580.6, 581.6, 582.6, 583.6, 584.6, 585.6, 586.6, 587.6, 588.6, 589.6, 590.6, 591.6, 592.6, 593.6, 594.6, 595.6, 596.6, 597.6, 598.6, 599.6, 600.6, 601.6, 602.6, 603.6, 604.6, 605.6, 606.6, 607.6, 608.6, 609.6, 610.6, 611.6, 612.6, 613.6, 614.6, 615.6, 616.6, 617.6, 618.6, 619.6, 620.6, 621.6, 622.6, 623.6, 624.6, 625.6, 626.6, 627.6, 628.6, 629.6, 630.6, 631.6, 632.6, 633.6, 634.6, 635.6, 636.6, 637.6, 638.6, 639.6, 640.6, 641.6, 642.6, 643.6, 644.6, 645.6, 646.6, 647.6, 648.6, 649.6, 650.6, 651.6, 652.6, 653.6, 654.6, 655.6, 656.6, 657.6, 658.6, 659.6, 660.7, 661.7, 662.7, 663.7, 664.7, 665.7, 666.7, 667.7, 668.7, 669.7, 670.7, 671.7, 672.7, 673.7, 674.7, 675.7, 676.7, 677.7, 678.7, 679.7, 680.7, 681.7, 682.7, 683.7, 684.7, 685.7, 686.7, 687.7, 688.7, 689.7, 690.7, 691.7, 692.7, 693.7, 694.7, 695.7, 696.7, 697.7, 698.7, 699.7, 700.7, 701.7, 702.7, 703.7, 704.7, 705.7, 706.7, 707.7, 708.7, 709.7, 710.7, 711.7, 712.7, 713.7, 714.7, 715.7, 716.7, 717.7, 718.7, 719.7, 720.7, 721.7, 722.7, 723.7, 724.7, 725.7, 726.7, 727.7, 728.7, 729.7, 730.7, 731.7, 732.7, 733.7, 734.7, 735.7, 736.7, 737.7, 738.7, 739.7, 740.7, 741.7, 742.7, 743.7, 744.7, 745.7, 746.7, 747.7, 748.7, 749.7, 750.7, 751.7, 752.7, 753.7, 754.7, 755.7, 756.7, 757.7, 758.7, 759.7, 760.7, 761.7, 762.8, 763.8, 764.8, 765.8, 766.8, 767.8, 768.8, 769.8, 770.8, 771.8, 772.8, 773.8, 774.8, 775.8, 776.8, 777.8, 778.8, 779.8, 780.8, 781.8, 782.8, 783.8, 784.8, 785.8, 786.8, 787.8, 788.8, 789.8, 790.8, 791.8, 792.8, 793.8, 794.8, 795.8, 796.8, 797.8, 798.8, 799.8, 800.8, 801.8, 802.8, 803.8, 804.8, 805.8, 806.8, 807.8, 808.8, 809.8, 810.8, 811.8, 812.8, 813.8, 814.3, 815.3, 816.3, 817.3, 818.3, 819.3, 820.3, 821.3, 822.3, 823.3, 824.3, 825.3, 826.3, 827.3, 828.3, 829.3, 830.3, 831.3, 832.3, 833.3, 834.3, 835.3, 836.3, 837.3, 838.3, 839.3, 840.3, 841.3, 842.3, 843.3, 844.3, 845.3, 846.3, 847.3, 848.3, 849.3, 850.3, 851.3, 852.3, 853.3, 854.3, 855.3, 856.3, 857.3, 858.3, 859.3, 860.3, 861.3, 862.3, 863.3, 864.4, 865.4, 866.4, 867.4, 868.4, 869.4, 870.4, 871.4, 872.4, 873.4, 874.4, 875.4, 876.4, 877.4, 878.4, 879.4, 880.4, 881.4, 882.4, 883.4, 884.4, 885.4, 886.4, 887.4, 888.4, 889.4, 890.4, 891.4, 892.4, 893.4, 894.4, 895.4, 896.4, 897.4, 898.4, 899.4, 900.4, 901.4, 902.4, 903.4, 904.4, 905.4, 906.4, 907.4, 908.4, 909.4, 910.4, 911.4, 912.4, 913.4, 914.4, 915.4, 916.4, 917.4, 918.4, 919.4, 920.4, 921.4, 922.4, 923.4, 924.4, 925.4, 926.4, 927.4, 928.4, 929.4, 930.4, 931.4, 932.4, 933.4, 934.4, 935.4, 936.4, 937.4, 938.4, 939.4, 940.4, 941.4, 942.4, 943.4, 944.4, 945.4, 946.4, 947.4, 948.4, 949.4, 950.4, 951.4, 952.4, 953.4, 954.4, 955.4, 956.4, 957.4, 958.4, 959.4, 960.4, 961.4, 962.4, 963.4, 964.4, 965.4, 966.5, 967.5, 968.5, 969.5, 970.5, 971.5, 972.5, 973.5, 974.5, 975.5, 976.5, 977.5, 978.5, 979.5, 980.5, 981.5, 982.5, 983.5, 984.5, 985.5, 986.5, 987.5, 988.5, 989.5, 990.5, 991.5, 992.5, 993.5, 994.5, 995.5, 996.5, 997.5, 998.5, 999.5, 1000.5, 1001.5, 1002.5, 1003.5, 1004.5, 1005.5, 1006.5, 1007.0, 1008.0, 1009.0, 1010.0, 1011.0, 1012.0, 1013.0, 1014.0, 1015.0, 1016.0, 1017.0, 1018.0, 1019.0, 1020.0, 1021.0, 1022.0, 1023.0, 1024.0, 1025.0, 1026.0, 1027.0, 1028.0, 1029.0, 1030.0, 1031.0, 1032.0, 1033.0, 1034.0, 1035.0, 1036.0, 1037.0, 1038.0, 1039.0, 1040.0, 1041.0, 1042.0, 1043.0, 1044.0, 1045.0, 1046.0, 1047.0, 1048.0, 1049.0, 1050.0, 1051.0, 1052.0, 1053.0, 1054.0, 1055.0, 1056.0, 1057.0, 1058.0, 1059.0, 1060.0, 1061.0, 1062.0, 1063.0, 1064.0, 1065.0, 1066.0, 1067.0, 1068.0, 1069.0, 1070.0, 1071.0, 1072.0, 1073.0, 1074.0, 1075.0, 1076.0, 1077.0, 1078.0, 1079.1, 1080.1, 1081.1, 1082.1, 1083.1, 1084.1, 1085.1, 1086.1, 1087.1, 1088.1, 1089.1, 1090.1, 1091.1, 1092.1, 1093.1, 1094.1, 1095.1, 1096.1, 1097.1, 1098.1, 1099.1, 1099.6, 1100.6, 1101.6, 1102.6, 1103.6, 1104.6, 1105.6, 1106.6, 1107.6, 1108.6, 1109.6, 1110.6, 1111.6, 1112.6, 1113.6, 1114.6, 1115.6, 1116.6, 1117.6, 1118.6, 1119.6, 1120.6, 1121.6, 1122.6, 1123.6, 1124.6, 1125.6, 1126.6, 1127.6, 1128.6, 1129.6, 1130.6, 1131.6, 1132.6, 1133.6, 1134.6, 1135.6, 1136.6, 1137.6, 1138.6, 1139.6, 1140.6, 1141.6, 1142.6, 1143.6, 1144.6, 1145.6, 1146.6, 1147.6, 1148.6, 1149.6, 1150.6, 1151.6, 1152.6, 1153.6, 1154.6, 1155.6, 1156.6, 1157.6, 1158.6, 1159.6, 1160.6, 1161.6, 1162.6, 1163.6, 1164.6, 1165.6, 1166.6, 1167.6, 1168.6, 1169.6, 1170.6, 1171.6, 1172.6, 1173.6, 1174.6, 1175.6, 1176.6, 1177.6, 1178.6, 1179.6, 1180.6, 1181.2, 1182.2, 1183.2, 1184.2, 1185.2, 1186.2, 1187.2, 1188.2, 1189.2, 1190.2, 1191.2, 1192.2, 1193.2, 1194.2, 1195.2, 1196.2, 1197.2, 1198.2, 1199.2, 1200.2, 1201.2, 1202.2, 1203.2, 1204.2, 1205.2, 1206.2, 1207.2, 1208.2, 1209.2, 1210.2, 1211.2, 1212.2, 1213.2, 1214.2, 1215.2, 1216.2, 1217.2, 1218.2, 1219.2, 1220.2, 1221.2, 1222.2, 1223.2, 1224.2, 1225.2, 1226.2, 1227.2, 1228.2, 1229.2, 1230.2, 1231.2, 1232.2, 1233.2, 1234.2, 1235.2, 1236.2, 1237.2, 1238.2, 1239.2, 1240.2, 1241.2, 1242.2, 1243.2, 1244.2, 1245.2, 1246.2, 1247.2, 1248.2, 1249.2, 1250.2, 1251.2, 1252.2, 1253.2, 1254.2, 1255.2, 1256.2, 1257.2, 1258.2, 1259.2, 1260.2, 1261.2, 1262.2, 1262.7, 1263.7, 1264.7, 1265.7, 1266.7, 1267.7, 1268.7, 1269.7, 1270.7, 1271.7, 1272.8, 1273.8, 1274.8, 1275.8, 1276.8, 1277.8, 1278.8, 1279.8, 1280.8, 1281.8, 1282.8, 1283.8, 1284.8, 1285.8, 1286.8, 1287.8, 1288.8, 1289.8, 1290.8, 1291.8, 1292.8, 1293.8, 1294.8, 1295.8, 1296.8, 1297.8, 1298.8, 1299.8, 1300.8, 1301.8, 1302.8, 1303.8, 1304.8, 1305.8, 1306.8, 1307.8, 1308.8, 1309.8, 1310.8, 1311.8, 1312.8, 1313.8, 1314.8, 1315.8, 1316.8, 1317.8, 1318.8, 1319.8, 1320.8, 1321.8, 1322.8, 1323.3, 1324.3, 1325.3, 1326.3, 1327.3, 1328.3, 1329.3, 1330.3, 1331.3, 1332.3, 1333.3, 1334.3, 1335.3, 1336.3, 1337.3, 1338.3, 1339.3, 1340.3, 1341.3, 1342.3, 1343.3, 1344.3, 1345.3, 1346.3, 1347.3, 1348.3, 1349.3, 1350.3, 1351.3, 1352.3, 1353.3, 1354.3, 1355.3, 1356.3, 1357.3, 1358.3, 1359.3, 1360.3, 1361.3, 1362.3, 1363.3, 1364.3, 1364.8, 1365.8, 1366.8, 1367.8, 1368.8, 1369.8, 1370.8, 1371.8, 1372.8, 1373.8, 1374.9, 1375.9, 1376.9, 1377.9, 1378.9, 1379.9, 1380.9, 1381.9, 1382.9, 1383.9, 1384.9, 1385.9, 1386.9, 1387.9, 1388.9, 1389.9, 1390.9, 1391.9, 1392.9, 1393.9, 1394.9, 1395.9, 1396.9, 1397.9, 1398.9, 1399.9, 1400.9, 1401.9, 1402.9, 1403.9, 1404.9, 1405.9, 1406.9, 1407.9, 1408.9, 1409.9, 1410.9, 1411.9, 1412.9, 1413.9, 1414.9, 1415.9, 1416.9, 1417.9, 1418.9, 1419.9, 1420.9, 1421.9, 1422.9, 1423.9, 1424.9, 1425.9, 1426.9, 1427.9, 1428.9, 1429.9, 1430.9, 1431.9, 1432.9, 1433.9, 1434.9, 1435.9, 1436.9, 1437.9, 1438.9, 1439.9, 1440.9, 1441.9, 1442.9, 1443.9, 1444.9, 1445.9, 1446.9, 1447.9, 1448.9, 1449.9, 1450.9, 1451.9, 1452.9, 1453.9, 1454.9, 1455.9, 1456.9, 1457.9, 1458.9, 1459.9, 1460.9, 1461.9, 1462.9, 1463.9, 1464.9, 1465.9, 1466.4, 1467.4, 1468.4, 1469.4, 1470.4, 1471.4, 1472.4, 1473.4, 1474.4, 1475.4, 1476.5, 1477.5, 1478.5, 1479.5, 1480.5, 1481.5, 1482.5, 1483.5, 1484.5, 1485.5, 1486.5, 1487.5, 1488.5, 1489.5, 1490.5, 1491.5, 1492.5, 1493.5, 1494.5, 1495.5, 1496.5, 1497.5, 1498.5, 1499.5, 1500.5, 1501.5, 1502.5, 1503.5, 1504.5, 1505.5, 1506.5, 1507.5, 1508.5, 1509.5, 1510.5, 1511.5, 1512.5, 1513.5, 1514.5, 1515.5, 1516.5, 1517.5, 1518.5, 1519.5, 1520.5, 1521.5, 1522.5, 1523.5, 1524.5, 1525.5, 1526.5, 1527.5, 1528.5, 1529.5, 1530.5, 1531.5, 1532.5, 1533.5, 1534.5, 1535.5, 1536.5, 1537.5, 1538.5, 1539.5, 1540.5, 1541.5, 1542.5, 1543.5, 1544.5, 1545.5, 1546.5, 1547.5, 1548.0, 1549.0, 1550.0, 1551.0, 1552.0, 1553.0, 1554.0, 1555.0, 1556.0, 1557.0, 1558.0, 1559.0, 1560.0, 1561.0, 1562.0, 1563.0, 1564.0, 1565.0, 1566.0, 1567.0, 1568.0, 1569.0, 1570.0, 1571.0, 1572.0, 1573.0, 1574.0, 1575.0, 1576.0, 1577.0, 1578.0, 1579.0, 1580.0, 1581.0, 1582.0, 1583.0, 1584.0, 1585.0, 1586.0, 1587.0, 1588.0, 1589.1, 1590.1, 1591.1, 1592.1, 1593.1, 1594.1, 1595.1, 1596.1, 1597.1, 1598.1, 1599.1, 1600.1, 1601.1, 1602.1, 1603.1, 1604.1, 1605.1, 1606.1, 1607.1, 1608.1, 1609.1, 1610.1, 1611.1, 1612.1, 1613.1, 1614.1, 1615.1, 1616.1, 1617.1, 1618.1, 1619.1, 1620.1, 1621.1, 1622.1, 1623.1, 1624.1, 1625.1, 1626.1, 1627.1, 1628.1, 1629.1, 1630.1, 1631.1, 1632.1, 1633.1, 1634.1, 1635.1, 1636.1, 1637.1, 1638.1, 1639.1, 1640.1, 1641.1, 1642.1, 1643.1, 1644.1, 1645.1, 1646.1, 1647.1, 1648.1, 1649.1, 1650.1, 1651.1, 1652.1, 1653.1, 1654.1, 1655.1, 1656.1, 1657.1, 1658.1, 1659.1, 1660.1, 1661.1, 1662.1, 1663.1, 1664.1, 1665.1, 1666.1, 1667.1, 1668.1, 1669.1, 1670.1, 1671.1, 1672.1, 1673.1, 1674.1, 1675.1, 1676.1, 1677.1, 1678.1, 1679.1, 1680.1, 1681.1, 1682.1, 1683.1, 1684.1, 1685.1, 1686.1, 1687.1, 1688.1, 1689.1, 1690.1, 1691.2, 1692.2, 1693.2, 1694.2, 1695.2, 1696.2, 1697.2, 1698.2, 1699.2, 1700.2, 1701.2, 1702.2, 1703.2, 1704.2, 1705.2, 1706.2, 1707.2, 1708.2, 1709.2, 1710.2, 1711.2, 1712.2, 1713.2, 1714.2, 1715.2, 1716.2, 1717.2, 1718.2, 1719.2, 1720.2, 1721.2, 1722.2, 1723.2, 1724.2, 1725.2, 1726.2, 1727.2, 1728.2, 1729.2, 1730.2, 1731.2, 1732.2, 1733.2, 1734.2, 1735.2, 1736.2, 1737.2, 1738.2, 1739.2, 1740.2, 1741.2, 1742.2, 1743.2, 1744.2, 1745.2, 1746.2, 1747.2, 1748.2, 1749.2, 1750.2, 1751.2, 1752.2, 1753.2, 1754.2, 1755.2, 1756.2, 1757.2, 1758.2, 1759.2, 1760.2, 1761.2, 1762.2, 1763.2, 1763.7, 1764.7, 1765.7, 1766.7, 1767.7, 1768.7, 1769.7, 1770.7, 1771.7, 1772.7, 1773.2, 1774.2, 1775.2, 1776.2, 1777.2, 1778.2, 1779.2, 1780.2, 1781.2, 1782.2, 1783.3, 1784.3, 1785.3, 1786.3, 1787.3, 1788.3, 1789.3, 1790.3, 1791.3, 1792.3, 1793.3, 1794.3, 1795.3, 1796.3, 1797.3, 1798.3, 1799.3, 1800.3, 1801.3, 1802.3, 1802.8, 1803.8, 1804.8, 1805.8, 1806.8, 1807.8, 1808.8, 1809.8, 1810.8, 1811.8, 1812.8, 1813.3, 1814.3, 1815.3, 1816.3, 1817.3, 1818.3, 1819.3, 1820.3, 1821.3, 1822.3, 1823.3, 1823.8, 1824.8, 1825.8, 1826.8, 1827.8, 1828.8, 1829.8, 1830.8, 1831.8, 1832.8, 1833.8, 1834.8, 1835.8, 1836.8, 1837.8, 1838.8, 1839.8, 1840.8, 1841.8, 1842.8, 1843.8, 1844.8, 1845.8, 1846.8, 1847.8, 1848.8, 1849.8, 1850.8, 1851.8, 1852.8, 1853.8, 1854.8, 1855.8, 1856.8, 1857.8, 1858.8, 1859.8, 1860.8, 1861.8, 1862.8, 1863.8, 1864.8, 1865.3, 1866.3, 1867.3, 1868.3, 1869.3, 1870.3, 1871.3, 1872.3, 1873.3, 1874.3, 1874.8, 1875.8, 1876.8, 1877.8, 1878.8, 1879.8, 1880.8, 1881.8, 1882.8, 1883.8, 1884.8, 1885.3, 1886.3, 1887.3, 1888.3, 1889.3, 1890.3, 1891.3, 1892.3, 1893.3, 1893.8, 1894.8, 1895.4, 1896.4, 1897.4, 1898.4, 1899.4, 1900.4, 1901.4, 1902.4, 1903.4, 1904.4, 1905.4, 1906.4, 1907.4, 1908.4, 1909.4, 1910.4, 1911.4, 1912.4, 1913.4, 1914.4, 1915.4, 1916.4, 1917.4, 1918.4, 1919.4, 1920.4, 1921.4, 1922.4, 1923.4, 1924.4, 1925.4, 1925.9, 1926.9, 1927.9, 1928.9, 1929.9, 1930.9, 1931.9, 1932.9, 1933.9, 1934.9, 1935.9, 1936.9, 1937.9, 1938.9, 1939.9, 1940.9, 1941.9, 1942.9, 1943.9, 1944.9, 1945.9, 1946.9, 1947.9, 1948.9, 1949.9, 1950.9, 1951.9, 1952.9, 1953.9, 1954.9, 1955.9, 1956.9, 1957.9, 1958.9, 1959.9, 1960.9, 1961.9, 1962.9, 1963.9, 1964.9, 1965.9, 1966.4, 1967.4, 1968.4, 1969.4, 1970.4, 1971.4, 1972.4, 1973.4, 1974.4, 1975.4, 1976.4, 1977.4, 1978.4, 1979.4, 1980.4, 1981.4, 1982.4, 1983.4, 1984.4, 1985.4, 1986.5, 1987.5, 1988.5, 1989.5, 1990.5, 1991.5, 1992.5, 1993.5, 1994.5, 1995.5, 1996.5, 1997.5, 1998.5, 1999.5, 2000.5, 2001.5, 2002.5, 2003.5, 2004.5, 2005.5, 2006.5, 2007.5, 2008.0, 2009.0, 2010.0, 2011.0, 2012.0, 2013.0, 2014.0, 2015.0, 2016.0, 2017.0, 2018.0, 2019.0, 2020.0, 2021.0, 2022.0, 2023.0, 2024.0, 2025.0, 2026.0, 2027.0, 2028.0, 2029.0, 2030.0, 2031.0, 2032.0, 2033.0, 2034.0, 2035.0, 2036.0, 2037.0, 2038.0, 2039.0, 2040.0, 2041.0, 2042.0, 2043.0, 2044.0, 2045.0, 2046.0, 2047.0, 2048.0, 2049.0, 2049.5, 2050.5, 2051.5, 2052.5, 2053.5, 2054.5, 2055.5, 2056.5, 2057.5, 2058.5, 2059.5, 2060.5, 2061.5, 2062.5, 2063.5, 2064.5, 2065.5, 2066.5, 2067.5, 2068.5, 2069.5, 2070.5, 2071.5, 2072.5, 2073.5, 2074.5, 2075.5, 2076.5, 2077.5, 2078.5, 2079.5, 2080.5, 2081.5, 2082.5, 2083.5, 2084.5, 2085.5, 2086.5, 2087.5, 2088.6, 2089.6, 2090.6, 2091.6, 2092.6, 2093.6, 2094.6, 2095.6, 2096.6, 2097.6, 2098.6, 2099.6, 2100.1, 2101.1, 2102.1, 2103.1, 2104.1, 2105.1, 2106.1, 2107.1, 2108.1, 2109.1, 2110.1, 2111.1, 2112.1, 2113.1, 2114.1, 2115.1, 2116.1, 2117.1, 2118.1, 2119.1, 2120.1, 2121.1, 2122.1, 2123.1, 2124.1, 2125.1, 2126.1, 2127.1, 2128.1, 2129.1, 2130.1, 2131.1, 2132.1, 2133.1, 2134.1, 2135.1, 2136.1, 2137.1, 2138.1, 2139.1, 2140.1, 2141.1, 2142.1, 2143.1, 2144.1, 2145.1, 2146.1, 2147.1, 2148.1, 2149.1, 2150.1, 2150.6, 2151.6, 2152.6, 2153.6, 2154.6, 2155.6, 2156.6, 2157.6, 2158.6, 2159.6, 2160.6, 2161.6, 2162.6, 2163.6, 2164.6, 2165.6, 2166.6, 2167.6, 2168.6, 2169.6, 2170.6, 2171.1, 2172.1, 2173.1, 2174.1, 2175.1, 2176.1, 2177.1, 2178.1, 2179.1, 2180.1, 2181.1, 2182.1, 2183.1, 2184.1, 2185.1, 2186.1, 2187.1, 2188.1, 2189.1, 2190.1, 2191.1, 2192.1, 2193.1, 2194.1, 2195.1, 2196.1, 2197.1, 2198.1, 2199.1, 2200.1, 2201.2, 2202.2, 2203.2, 2204.2, 2205.2, 2206.2, 2207.2, 2208.2, 2209.2, 2210.2, 2211.2, 2212.2, 2213.2, 2214.2, 2215.2, 2216.2, 2217.2, 2218.2, 2219.2, 2220.2, 2221.2, 2222.2, 2222.7, 2223.7, 2224.7, 2225.7, 2226.7, 2227.7, 2228.7, 2229.7, 2230.7, 2231.7, 2232.7, 2233.7, 2234.7, 2235.7, 2236.7, 2237.7, 2238.7, 2239.7, 2240.7, 2241.7, 2242.7, 2243.7, 2244.7, 2245.7, 2246.7, 2247.7, 2248.7, 2249.7, 2250.7, 2251.7, 2252.7, 2253.7, 2254.2, 2255.2, 2256.2, 2257.2, 2258.2, 2259.2, 2260.2, 2261.2, 2262.2, 2262.7, 2263.7, 2264.7, 2265.7, 2266.7, 2267.7, 2268.7, 2269.7, 2270.7, 2271.7, 2272.7, 2273.2, 2274.2, 2275.2, 2276.2, 2277.2, 2278.2, 2279.2, 2280.2, 2281.2, 2282.2, 2283.2, 2283.7, 2284.7, 2285.7, 2286.7, 2287.7, 2288.7, 2289.7, 2290.7, 2291.7, 2292.8, 2293.8, 2294.8, 2295.8, 2296.8, 2297.8, 2298.8, 2299.8, 2300.8, 2301.8, 2302.8, 2303.8, 2304.3, 2305.3, 2306.3, 2307.3, 2308.3, 2309.3, 2310.3, 2311.3, 2312.3, 2313.3, 2314.3, 2314.8, 2315.8, 2316.8, 2317.8, 2318.8, 2319.8, 2320.8, 2321.8, 2322.8, 2323.8, 2324.8, 2325.3, 2326.3, 2327.3, 2328.3, 2329.3, 2330.3, 2331.3, 2332.3, 2333.3, 2334.3, 2334.8, 2335.8, 2336.8, 2337.8, 2338.8, 2339.8, 2340.8, 2341.8, 2342.8, 2343.8, 2344.8, 2345.8, 2346.8, 2347.8, 2348.8, 2349.8, 2350.8, 2351.8, 2352.8, 2353.8, 2354.8, 2355.3, 2356.3, 2357.3, 2358.3, 2359.3, 2360.3, 2361.3, 2362.3, 2363.3, 2364.3, 2365.3, 2366.3, 2367.3, 2368.3, 2369.3, 2370.3, 2371.3, 2372.3, 2373.3, 2374.3, 2375.3, 2376.3, 2377.3, 2378.3, 2379.3, 2380.3, 2381.3, 2382.3, 2383.3, 2384.3, 2385.3, 2385.8, 2386.8, 2387.8, 2388.8, 2389.8, 2390.8, 2391.8, 2392.8, 2393.8, 2394.8, 2395.3, 2396.3, 2397.3, 2398.3, 2399.3, 2400.3, 2401.3, 2402.3, 2403.3, 2404.3, 2405.4, 2406.4, 2407.4, 2408.4, 2409.4, 2410.4, 2411.4, 2412.4, 2413.4, 2414.4, 2415.4, 2415.9, 2416.9, 2417.9, 2418.9, 2419.9, 2420.9, 2421.9, 2422.9, 2423.9, 2424.9, 2425.9, 2426.4, 2427.4, 2428.4, 2429.4, 2430.4, 2431.4, 2432.4, 2433.4, 2434.4, 2435.4, 2436.4, 2436.9, 2437.9, 2438.9, 2439.9, 2440.9, 2441.9, 2442.9, 2443.9, 2444.9, 2445.9, 2446.9, 2447.4, 2448.4, 2449.4, 2450.4, 2451.4, 2452.4, 2453.4, 2454.4, 2455.4, 2456.4, 2457.4, 2457.9, 2458.9, 2459.9, 2460.9, 2461.9, 2462.9, 2463.9, 2464.9, 2465.9, 2466.9, 2467.9, 2468.9, 2469.9, 2470.9, 2471.9, 2472.9, 2473.9, 2474.9, 2475.9, 2476.9, 2477.9, 2478.9, 2479.9, 2480.9, 2481.9, 2482.9, 2483.9, 2484.9, 2485.9, 2486.9, 2487.9, 2488.4, 2489.4, 2490.4, 2491.4, 2492.4, 2493.4, 2494.4, 2495.4, 2496.4, 2497.5, 2498.5, 2499.5, 2500.5, 2501.5, 2502.5, 2503.5, 2504.5, 2505.5, 2506.5, 2507.5, 2508.0, 2509.0, 2510.0, 2511.0, 2512.0, 2513.0, 2514.0, 2515.0, 2516.0, 2517.0, 2518.0, 2519.0, 2520.0, 2521.0, 2522.0, 2523.0, 2524.0, 2525.0, 2526.0, 2527.0, 2528.0, 2528.5, 2529.5, 2530.5, 2531.5, 2532.5, 2533.5, 2534.5, 2535.5, 2536.5, 2537.5, 2538.0, 2539.0, 2540.0, 2541.0, 2542.0, 2543.0, 2544.0, 2545.0, 2546.0, 2547.0, 2548.0, 2549.0, 2549.5, 2550.5, 2551.5, 2552.5, 2553.5, 2554.5, 2555.5, 2556.5, 2557.5, 2558.5, 2559.5, 2560.5, 2561.5, 2562.5, 2563.5, 2564.5, 2565.5, 2566.5, 2567.5, 2568.5, 2569.0, 2570.0, 2571.0, 2572.0, 2573.0, 2574.0, 2575.0, 2576.0, 2577.0, 2578.0, 2579.0, 2580.0, 2580.5, 2581.5, 2582.5, 2583.5, 2584.5, 2585.5, 2586.5, 2587.5, 2588.5, 2589.5, 2590.5, 2591.5, 2592.5, 2593.5, 2594.5, 2595.5, 2596.5, 2597.5, 2598.5, 2599.5, 2600.1, 2601.1, 2602.1, 2603.1, 2604.1, 2605.1, 2606.1, 2607.1, 2608.1, 2609.1, 2609.6, 2610.6, 2611.6, 2612.6, 2613.6, 2614.6, 2615.6, 2616.6, 2617.6, 2618.6, 2619.6, 2620.6, 2621.6, 2622.6, 2623.6, 2624.6, 2625.6, 2626.6, 2627.6, 2628.6, 2629.6, 2630.1, 2631.1, 2632.1, 2633.1, 2634.1, 2635.1, 2636.1, 2637.1, 2638.1, 2639.1, 2640.1, 2641.1, 2642.1, 2643.1, 2644.1, 2645.1, 2646.1, 2647.1, 2648.1, 2649.1, 2650.1, 2651.1, 2652.1, 2653.1, 2654.1, 2655.1, 2656.1, 2657.1, 2658.1, 2659.1, 2660.1, 2661.1, 2662.1, 2662.6, 2663.6, 2664.6, 2665.6, 2666.6}
time =
  {9.62347748E8, 9.62347749E8, 9.6234775E8, 9.62347751E8, 9.62347752E8, 9.62347753E8, 9.62347754E8, 9.62347755E8, 9.62347756E8, 9.62347757E8, 9.62347758E8, 9.62347759E8, 9.6234776E8, 9.62347761E8, 9.62347762E8, 9.62347763E8, 9.62347764E8, 9.62347765E8, 9.62347766E8, 9.62347767E8, 9.62347768E8, 9.62347769E8, 9.6234777E8, 9.62347771E8, 9.62347772E8, 9.62347773E8, 9.62347774E8, 9.62347775E8, 9.62347776E8, 9.62347777E8, 9.62347778E8, 9.62347779E8, 9.6234778E8, 9.62347781E8, 9.62347782E8, 9.62347783E8, 9.62347784E8, 9.62347785E8, 9.62347786E8, 9.62347787E8, 9.62347788E8, 9.62347789E8, 9.6234779E8, 9.62347791E8, 9.62347792E8, 9.62347793E8, 9.62347794E8, 9.62347795E8, 9.62347796E8, 9.62347797E8, 9.62347798E8, 9.62347799E8, 9.623478E8, 9.62347801E8, 9.62347802E8, 9.62347803E8, 9.62347804E8, 9.62347805E8, 9.62347806E8, 9.62347807E8, 9.623478081E8, 9.623478091E8, 9.623478101E8, 9.623478111E8, 9.623478121E8, 9.623478131E8, 9.623478141E8, 9.623478151E8, 9.623478161E8, 9.623478171E8, 9.623478181E8, 9.623478191E8, 9.623478201E8, 9.623478211E8, 9.623478221E8, 9.623478231E8, 9.623478241E8, 9.623478251E8, 9.623478261E8, 9.623478271E8, 9.623478281E8, 9.623478291E8, 9.623478301E8, 9.623478311E8, 9.623478321E8, 9.623478331E8, 9.623478341E8, 9.623478351E8, 9.623478361E8, 9.623478371E8, 9.623478381E8, 9.623478391E8, 9.623478401E8, 9.623478411E8, 9.623478421E8, 9.623478431E8, 9.623478441E8, 9.623478451E8, 9.623478461E8, 9.623478471E8, 9.623478481E8, 9.623478491E8, 9.623478501E8, 9.623478511E8, 9.623478521E8, 9.623478531E8, 9.623478541E8, 9.623478551E8, 9.623478561E8, 9.623478571E8, 9.623478581E8, 9.623478591E8, 9.623478601E8, 9.623478611E8, 9.623478621E8, 9.623478631E8, 9.623478641E8, 9.623478651E8, 9.623478661E8, 9.623478671E8, 9.623478681E8, 9.623478691E8, 9.623478701E8, 9.623478711E8, 9.623478721E8, 9.623478731E8, 9.623478741E8, 9.623478751E8, 9.623478761E8, 9.623478771E8, 9.623478781E8, 9.623478791E8, 9.623478801E8, 9.623478811E8, 9.623478821E8, 9.623478831E8, 9.623478841E8, 9.623478851E8, 9.623478861E8, 9.623478871E8, 9.623478881E8, 9.623478891E8, 9.623478901E8, 9.623478911E8, 9.623478921E8, 9.623478931E8, 9.623478941E8, 9.623478951E8, 9.623478961E8, 9.623478971E8, 9.623478981E8, 9.623478991E8, 9.623479001E8, 9.623479011E8, 9.623479021E8, 9.623479031E8, 9.623479041E8, 9.623479051E8, 9.623479061E8, 9.623479072E8, 9.623479082E8, 9.623479092E8, 9.623479102E8, 9.623479112E8, 9.623479122E8, 9.623479132E8, 9.623479142E8, 9.623479152E8, 9.623479162E8, 9.623479172E8, 9.623479182E8, 9.623479192E8, 9.623479202E8, 9.623479212E8, 9.623479222E8, 9.623479232E8, 9.623479242E8, 9.623479252E8, 9.623479262E8, 9.623479272E8, 9.623479282E8, 9.623479292E8, 9.623479302E8, 9.623479312E8, 9.623479322E8, 9.623479332E8, 9.623479342E8, 9.623479352E8, 9.623479362E8, 9.623479372E8, 9.623479382E8, 9.623479392E8, 9.623479402E8, 9.623479412E8, 9.623479422E8, 9.623479432E8, 9.623479442E8, 9.623479452E8, 9.623479462E8, 9.623479472E8, 9.623479482E8, 9.623479492E8, 9.623479502E8, 9.623479512E8, 9.623479522E8, 9.623479532E8, 9.623479542E8, 9.623479552E8, 9.623479562E8, 9.623479572E8, 9.623479582E8, 9.623479592E8, 9.623479602E8, 9.623479612E8, 9.623479622E8, 9.623479632E8, 9.623479642E8, 9.623479652E8, 9.623479662E8, 9.623479672E8, 9.623479682E8, 9.623479692E8, 9.623479702E8, 9.623479712E8, 9.623479722E8, 9.623479732E8, 9.623479742E8, 9.623479752E8, 9.623479762E8, 9.623479772E8, 9.623479782E8, 9.623479792E8, 9.623479802E8, 9.623479812E8, 9.623479822E8, 9.623479832E8, 9.623479842E8, 9.623479852E8, 9.623479862E8, 9.623479872E8, 9.623479882E8, 9.623479892E8, 9.623479902E8, 9.623479912E8, 9.623479922E8, 9.623479932E8, 9.623479942E8, 9.623479952E8, 9.623479962E8, 9.623479972E8, 9.623479982E8, 9.623479992E8, 9.623480002E8, 9.623480012E8, 9.623480022E8, 9.623480032E8, 9.623480042E8, 9.623480052E8, 9.623480062E8, 9.623480072E8, 9.623480082E8, 9.623480092E8, 9.623480102E8, 9.623480113E8, 9.623480123E8, 9.623480133E8, 9.623480143E8, 9.623480153E8, 9.623480163E8, 9.623480173E8, 9.623480183E8, 9.623480193E8, 9.623480203E8, 9.623480213E8, 9.623480223E8, 9.623480233E8, 9.623480243E8, 9.623480253E8, 9.623480263E8, 9.623480273E8, 9.623480283E8, 9.623480293E8, 9.623480303E8, 9.623480313E8, 9.623480323E8, 9.623480333E8, 9.623480343E8, 9.623480353E8, 9.623480363E8, 9.623480373E8, 9.623480383E8, 9.623480393E8, 9.623480403E8, 9.623480413E8, 9.623480423E8, 9.623480433E8, 9.623480443E8, 9.623480453E8, 9.623480463E8, 9.623480473E8, 9.623480483E8, 9.623480493E8, 9.623480503E8, 9.623480513E8, 9.623480523E8, 9.623480533E8, 9.623480543E8, 9.623480553E8, 9.623480563E8, 9.623480573E8, 9.623480583E8, 9.623480593E8, 9.623480603E8, 9.623480613E8, 9.623480623E8, 9.623480633E8, 9.623480643E8, 9.623480653E8, 9.623480663E8, 9.623480673E8, 9.623480683E8, 9.623480693E8, 9.623480703E8, 9.623480713E8, 9.623480723E8, 9.623480733E8, 9.623480743E8, 9.623480753E8, 9.623480763E8, 9.623480773E8, 9.623480783E8, 9.623480793E8, 9.623480803E8, 9.623480813E8, 9.623480823E8, 9.623480833E8, 9.623480843E8, 9.623480853E8, 9.623480863E8, 9.623480873E8, 9.623480883E8, 9.623480893E8, 9.623480903E8, 9.623480913E8, 9.623480923E8, 9.623480933E8, 9.623480943E8, 9.623480953E8, 9.623480963E8, 9.623480973E8, 9.623480983E8, 9.623480993E8, 9.623481003E8, 9.623481013E8, 9.623481023E8, 9.623481033E8, 9.623481043E8, 9.623481053E8, 9.623481063E8, 9.623481073E8, 9.623481083E8, 9.623481093E8, 9.623481103E8, 9.623481113E8, 9.623481123E8, 9.623481134E8, 9.623481144E8, 9.623481154E8, 9.623481164E8, 9.623481174E8, 9.623481184E8, 9.623481194E8, 9.623481204E8, 9.623481214E8, 9.623481224E8, 9.623481234E8, 9.623481244E8, 9.623481254E8, 9.623481264E8, 9.623481274E8, 9.623481284E8, 9.623481294E8, 9.623481304E8, 9.623481314E8, 9.623481324E8, 9.623481334E8, 9.623481344E8, 9.623481354E8, 9.623481364E8, 9.623481374E8, 9.623481384E8, 9.623481394E8, 9.623481404E8, 9.623481414E8, 9.623481424E8, 9.623481434E8, 9.623481444E8, 9.623481454E8, 9.623481464E8, 9.623481474E8, 9.623481484E8, 9.623481494E8, 9.623481504E8, 9.623481514E8, 9.623481524E8, 9.623481534E8, 9.623481544E8, 9.623481554E8, 9.623481564E8, 9.623481574E8, 9.623481584E8, 9.623481594E8, 9.623481604E8, 9.623481614E8, 9.623481624E8, 9.623481634E8, 9.623481644E8, 9.623481654E8, 9.623481664E8, 9.623481674E8, 9.623481684E8, 9.623481694E8, 9.623481704E8, 9.623481714E8, 9.623481724E8, 9.623481734E8, 9.623481744E8, 9.623481754E8, 9.623481764E8, 9.623481774E8, 9.623481784E8, 9.623481794E8, 9.623481804E8, 9.623481814E8, 9.623481824E8, 9.623481834E8, 9.623481844E8, 9.623481854E8, 9.623481864E8, 9.623481874E8, 9.623481884E8, 9.623481894E8, 9.623481904E8, 9.623481914E8, 9.623481924E8, 9.623481934E8, 9.623481944E8, 9.623481954E8, 9.623481964E8, 9.623481974E8, 9.623481984E8, 9.623481994E8, 9.623482004E8, 9.623482014E8, 9.623482024E8, 9.623482034E8, 9.623482044E8, 9.623482055E8, 9.623482065E8, 9.623482075E8, 9.623482085E8, 9.623482095E8, 9.623482105E8, 9.623482115E8, 9.623482125E8, 9.623482135E8, 9.623482145E8, 9.623482155E8, 9.623482165E8, 9.623482175E8, 9.623482185E8, 9.623482195E8, 9.623482205E8, 9.623482215E8, 9.623482225E8, 9.623482235E8, 9.623482245E8, 9.623482255E8, 9.623482265E8, 9.623482275E8, 9.623482285E8, 9.623482295E8, 9.623482305E8, 9.623482315E8, 9.623482325E8, 9.623482335E8, 9.623482345E8, 9.623482355E8, 9.623482365E8, 9.623482375E8, 9.623482385E8, 9.623482395E8, 9.623482405E8, 9.623482415E8, 9.623482425E8, 9.623482435E8, 9.623482445E8, 9.623482455E8, 9.623482465E8, 9.623482475E8, 9.623482485E8, 9.623482495E8, 9.623482505E8, 9.623482515E8, 9.623482525E8, 9.623482535E8, 9.623482545E8, 9.623482555E8, 9.623482565E8, 9.623482575E8, 9.623482585E8, 9.623482595E8, 9.623482605E8, 9.623482615E8, 9.623482625E8, 9.623482635E8, 9.623482645E8, 9.623482655E8, 9.623482665E8, 9.623482675E8, 9.623482685E8, 9.623482695E8, 9.623482705E8, 9.623482715E8, 9.623482725E8, 9.623482735E8, 9.623482745E8, 9.623482755E8, 9.623482765E8, 9.623482775E8, 9.623482785E8, 9.623482795E8, 9.623482805E8, 9.623482815E8, 9.623482825E8, 9.623482835E8, 9.623482845E8, 9.623482855E8, 9.623482865E8, 9.623482875E8, 9.623482885E8, 9.623482895E8, 9.623482905E8, 9.623482915E8, 9.623482925E8, 9.623482935E8, 9.623482945E8, 9.623482955E8, 9.623482965E8, 9.623482975E8, 9.623482985E8, 9.623482995E8, 9.623483005E8, 9.623483015E8, 9.623483025E8, 9.623483035E8, 9.623483045E8, 9.623483055E8, 9.623483065E8, 9.623483075E8, 9.623483085E8, 9.623483095E8, 9.623483105E8, 9.623483115E8, 9.623483125E8, 9.623483135E8, 9.623483145E8, 9.623483155E8, 9.623483165E8, 9.623483176E8, 9.623483186E8, 9.623483196E8, 9.623483206E8, 9.623483216E8, 9.623483226E8, 9.623483236E8, 9.623483246E8, 9.623483256E8, 9.623483266E8, 9.623483276E8, 9.623483286E8, 9.623483296E8, 9.623483306E8, 9.623483316E8, 9.623483326E8, 9.623483336E8, 9.623483346E8, 9.623483356E8, 9.623483366E8, 9.623483376E8, 9.623483386E8, 9.623483396E8, 9.623483406E8, 9.623483416E8, 9.623483426E8, 9.623483436E8, 9.623483446E8, 9.623483456E8, 9.623483466E8, 9.623483476E8, 9.623483486E8, 9.623483496E8, 9.623483506E8, 9.623483516E8, 9.623483526E8, 9.623483536E8, 9.623483546E8, 9.623483556E8, 9.623483566E8, 9.623483576E8, 9.623483586E8, 9.623483596E8, 9.623483606E8, 9.623483616E8, 9.623483626E8, 9.623483636E8, 9.623483646E8, 9.623483656E8, 9.623483666E8, 9.623483676E8, 9.623483686E8, 9.623483696E8, 9.623483706E8, 9.623483716E8, 9.623483726E8, 9.623483736E8, 9.623483746E8, 9.623483756E8, 9.623483766E8, 9.623483776E8, 9.623483786E8, 9.623483796E8, 9.623483806E8, 9.623483816E8, 9.623483826E8, 9.623483836E8, 9.623483846E8, 9.623483856E8, 9.623483866E8, 9.623483876E8, 9.623483886E8, 9.623483896E8, 9.623483906E8, 9.623483916E8, 9.623483926E8, 9.623483936E8, 9.623483946E8, 9.623483956E8, 9.623483966E8, 9.623483976E8, 9.623483986E8, 9.623483996E8, 9.623484006E8, 9.623484016E8, 9.623484026E8, 9.623484036E8, 9.623484046E8, 9.623484056E8, 9.623484066E8, 9.623484076E8, 9.623484086E8, 9.623484097E8, 9.623484107E8, 9.623484117E8, 9.623484127E8, 9.623484137E8, 9.623484147E8, 9.623484157E8, 9.623484167E8, 9.623484177E8, 9.623484187E8, 9.623484197E8, 9.623484207E8, 9.623484217E8, 9.623484227E8, 9.623484237E8, 9.623484247E8, 9.623484257E8, 9.623484267E8, 9.623484277E8, 9.623484287E8, 9.623484297E8, 9.623484307E8, 9.623484317E8, 9.623484327E8, 9.623484337E8, 9.623484347E8, 9.623484357E8, 9.623484367E8, 9.623484377E8, 9.623484387E8, 9.623484397E8, 9.623484407E8, 9.623484417E8, 9.623484427E8, 9.623484437E8, 9.623484447E8, 9.623484457E8, 9.623484467E8, 9.623484477E8, 9.623484487E8, 9.623484497E8, 9.623484507E8, 9.623484517E8, 9.623484527E8, 9.623484537E8, 9.623484547E8, 9.623484557E8, 9.623484567E8, 9.623484577E8, 9.623484587E8, 9.623484597E8, 9.623484607E8, 9.623484617E8, 9.623484627E8, 9.623484637E8, 9.623484647E8, 9.623484657E8, 9.623484667E8, 9.623484677E8, 9.623484687E8, 9.623484697E8, 9.623484707E8, 9.623484717E8, 9.623484727E8, 9.623484737E8, 9.623484747E8, 9.623484757E8, 9.623484767E8, 9.623484777E8, 9.623484787E8, 9.623484797E8, 9.623484807E8, 9.623484817E8, 9.623484827E8, 9.623484837E8, 9.623484847E8, 9.623484857E8, 9.623484867E8, 9.623484877E8, 9.623484887E8, 9.623484897E8, 9.623484907E8, 9.623484917E8, 9.623484927E8, 9.623484937E8, 9.623484947E8, 9.623484957E8, 9.623484967E8, 9.623484977E8, 9.623484987E8, 9.623484997E8, 9.623485007E8, 9.623485017E8, 9.623485027E8, 9.623485037E8, 9.623485047E8, 9.623485057E8, 9.623485067E8, 9.623485077E8, 9.623485087E8, 9.623485097E8, 9.623485107E8, 9.623485118E8, 9.623485128E8, 9.623485138E8, 9.623485148E8, 9.623485158E8, 9.623485168E8, 9.623485178E8, 9.623485188E8, 9.623485198E8, 9.623485208E8, 9.623485218E8, 9.623485228E8, 9.623485238E8, 9.623485248E8, 9.623485258E8, 9.623485268E8, 9.623485278E8, 9.623485288E8, 9.623485298E8, 9.623485308E8, 9.623485318E8, 9.623485328E8, 9.623485338E8, 9.623485348E8, 9.623485358E8, 9.623485368E8, 9.623485378E8, 9.623485388E8, 9.623485398E8, 9.623485408E8, 9.623485418E8, 9.623485428E8, 9.623485438E8, 9.623485448E8, 9.623485458E8, 9.623485468E8, 9.623485478E8, 9.623485488E8, 9.623485498E8, 9.623485508E8, 9.623485518E8, 9.623485528E8, 9.623485538E8, 9.623485548E8, 9.623485558E8, 9.623485568E8, 9.623485578E8, 9.623485588E8, 9.623485598E8, 9.623485608E8, 9.623485618E8, 9.623485628E8, 9.623485633E8, 9.623485643E8, 9.623485653E8, 9.623485663E8, 9.623485673E8, 9.623485683E8, 9.623485693E8, 9.623485703E8, 9.623485713E8, 9.623485723E8, 9.623485733E8, 9.623485743E8, 9.623485753E8, 9.623485763E8, 9.623485773E8, 9.623485783E8, 9.623485793E8, 9.623485803E8, 9.623485813E8, 9.623485823E8, 9.623485833E8, 9.623485843E8, 9.623485853E8, 9.623485863E8, 9.623485873E8, 9.623485883E8, 9.623485893E8, 9.623485903E8, 9.623485913E8, 9.623485923E8, 9.623485933E8, 9.623485943E8, 9.623485953E8, 9.623485963E8, 9.623485973E8, 9.623485983E8, 9.623485993E8, 9.623486003E8, 9.623486013E8, 9.623486023E8, 9.623486033E8, 9.623486043E8, 9.623486053E8, 9.623486063E8, 9.623486073E8, 9.623486083E8, 9.623486093E8, 9.623486103E8, 9.623486113E8, 9.623486123E8, 9.623486134E8, 9.623486144E8, 9.623486154E8, 9.623486164E8, 9.623486174E8, 9.623486184E8, 9.623486194E8, 9.623486204E8, 9.623486214E8, 9.623486224E8, 9.623486234E8, 9.623486244E8, 9.623486254E8, 9.623486264E8, 9.623486274E8, 9.623486284E8, 9.623486294E8, 9.623486304E8, 9.623486314E8, 9.623486324E8, 9.623486334E8, 9.623486344E8, 9.623486354E8, 9.623486364E8, 9.623486374E8, 9.623486384E8, 9.623486394E8, 9.623486404E8, 9.623486414E8, 9.623486424E8, 9.623486434E8, 9.623486444E8, 9.623486454E8, 9.623486464E8, 9.623486474E8, 9.623486484E8, 9.623486494E8, 9.623486504E8, 9.623486514E8, 9.623486524E8, 9.623486534E8, 9.623486544E8, 9.623486554E8, 9.623486564E8, 9.623486574E8, 9.623486584E8, 9.623486594E8, 9.623486604E8, 9.623486614E8, 9.623486624E8, 9.623486634E8, 9.623486644E8, 9.623486654E8, 9.623486664E8, 9.623486674E8, 9.623486684E8, 9.623486694E8, 9.623486704E8, 9.623486714E8, 9.623486724E8, 9.623486734E8, 9.623486744E8, 9.623486754E8, 9.623486764E8, 9.623486774E8, 9.623486784E8, 9.623486794E8, 9.623486804E8, 9.623486814E8, 9.623486824E8, 9.623486834E8, 9.623486844E8, 9.623486854E8, 9.623486864E8, 9.623486874E8, 9.623486884E8, 9.623486894E8, 9.623486904E8, 9.623486914E8, 9.623486924E8, 9.623486934E8, 9.623486944E8, 9.623486954E8, 9.623486964E8, 9.623486974E8, 9.623486984E8, 9.623486994E8, 9.623487004E8, 9.623487014E8, 9.623487024E8, 9.623487034E8, 9.623487044E8, 9.623487054E8, 9.623487064E8, 9.623487074E8, 9.623487084E8, 9.623487094E8, 9.623487104E8, 9.623487114E8, 9.623487124E8, 9.623487134E8, 9.623487144E8, 9.623487155E8, 9.623487165E8, 9.623487175E8, 9.623487185E8, 9.623487195E8, 9.623487205E8, 9.623487215E8, 9.623487225E8, 9.623487235E8, 9.623487245E8, 9.623487255E8, 9.623487265E8, 9.623487275E8, 9.623487285E8, 9.623487295E8, 9.623487305E8, 9.623487315E8, 9.623487325E8, 9.623487335E8, 9.623487345E8, 9.623487355E8, 9.623487365E8, 9.623487375E8, 9.623487385E8, 9.623487395E8, 9.623487405E8, 9.623487415E8, 9.623487425E8, 9.623487435E8, 9.623487445E8, 9.623487455E8, 9.623487465E8, 9.623487475E8, 9.623487485E8, 9.623487495E8, 9.623487505E8, 9.623487515E8, 9.623487525E8, 9.623487535E8, 9.623487545E8, 9.623487555E8, 9.62348756E8, 9.62348757E8, 9.62348758E8, 9.62348759E8, 9.6234876E8, 9.62348761E8, 9.62348762E8, 9.62348763E8, 9.62348764E8, 9.62348765E8, 9.62348766E8, 9.62348767E8, 9.62348768E8, 9.62348769E8, 9.6234877E8, 9.62348771E8, 9.62348772E8, 9.62348773E8, 9.62348774E8, 9.62348775E8, 9.62348776E8, 9.62348777E8, 9.62348778E8, 9.62348779E8, 9.6234878E8, 9.62348781E8, 9.62348782E8, 9.62348783E8, 9.62348784E8, 9.62348785E8, 9.62348786E8, 9.62348787E8, 9.62348788E8, 9.62348789E8, 9.6234879E8, 9.62348791E8, 9.62348792E8, 9.62348793E8, 9.62348794E8, 9.62348795E8, 9.62348796E8, 9.62348797E8, 9.62348798E8, 9.62348799E8, 9.623488E8, 9.62348801E8, 9.62348802E8, 9.62348803E8, 9.62348804E8, 9.62348805E8, 9.62348806E8, 9.62348807E8, 9.62348808E8, 9.62348809E8, 9.6234881E8, 9.62348811E8, 9.62348812E8, 9.62348813E8, 9.62348814E8, 9.62348815E8, 9.62348816E8, 9.62348817E8, 9.62348818E8, 9.62348819E8, 9.6234882E8, 9.62348821E8, 9.62348822E8, 9.62348823E8, 9.62348824E8, 9.62348825E8, 9.62348826E8, 9.62348827E8, 9.623488281E8, 9.623488291E8, 9.623488301E8, 9.623488311E8, 9.623488321E8, 9.623488331E8, 9.623488341E8, 9.623488351E8, 9.623488361E8, 9.623488371E8, 9.623488381E8, 9.623488391E8, 9.623488401E8, 9.623488411E8, 9.623488421E8, 9.623488431E8, 9.623488441E8, 9.623488451E8, 9.623488461E8, 9.623488471E8, 9.623488481E8, 9.623488486E8, 9.623488496E8, 9.623488506E8, 9.623488516E8, 9.623488526E8, 9.623488536E8, 9.623488546E8, 9.623488556E8, 9.623488566E8, 9.623488576E8, 9.623488586E8, 9.623488596E8, 9.623488606E8, 9.623488616E8, 9.623488626E8, 9.623488636E8, 9.623488646E8, 9.623488656E8, 9.623488666E8, 9.623488676E8, 9.623488686E8, 9.623488696E8, 9.623488706E8, 9.623488716E8, 9.623488726E8, 9.623488736E8, 9.623488746E8, 9.623488756E8, 9.623488766E8, 9.623488776E8, 9.623488786E8, 9.623488796E8, 9.623488806E8, 9.623488816E8, 9.623488826E8, 9.623488836E8, 9.623488846E8, 9.623488856E8, 9.623488866E8, 9.623488876E8, 9.623488886E8, 9.623488896E8, 9.623488906E8, 9.623488916E8, 9.623488926E8, 9.623488936E8, 9.623488946E8, 9.623488956E8, 9.623488966E8, 9.623488976E8, 9.623488986E8, 9.623488996E8, 9.623489006E8, 9.623489016E8, 9.623489026E8, 9.623489036E8, 9.623489046E8, 9.623489056E8, 9.623489066E8, 9.623489076E8, 9.623489086E8, 9.623489096E8, 9.623489106E8, 9.623489116E8, 9.623489126E8, 9.623489136E8, 9.623489146E8, 9.623489156E8, 9.623489166E8, 9.623489176E8, 9.623489186E8, 9.623489196E8, 9.623489206E8, 9.623489216E8, 9.623489226E8, 9.623489236E8, 9.623489246E8, 9.623489256E8, 9.623489266E8, 9.623489276E8, 9.623489286E8, 9.623489296E8, 9.623489302E8, 9.623489312E8, 9.623489322E8, 9.623489332E8, 9.623489342E8, 9.623489352E8, 9.623489362E8, 9.623489372E8, 9.623489382E8, 9.623489392E8, 9.623489402E8, 9.623489412E8, 9.623489422E8, 9.623489432E8, 9.623489442E8, 9.623489452E8, 9.623489462E8, 9.623489472E8, 9.623489482E8, 9.623489492E8, 9.623489502E8, 9.623489512E8, 9.623489522E8, 9.623489532E8, 9.623489542E8, 9.623489552E8, 9.623489562E8, 9.623489572E8, 9.623489582E8, 9.623489592E8, 9.623489602E8, 9.623489612E8, 9.623489622E8, 9.623489632E8, 9.623489642E8, 9.623489652E8, 9.623489662E8, 9.623489672E8, 9.623489682E8, 9.623489692E8, 9.623489702E8, 9.623489712E8, 9.623489722E8, 9.623489732E8, 9.623489742E8, 9.623489752E8, 9.623489762E8, 9.623489772E8, 9.623489782E8, 9.623489792E8, 9.623489802E8, 9.623489812E8, 9.623489822E8, 9.623489832E8, 9.623489842E8, 9.623489852E8, 9.623489862E8, 9.623489872E8, 9.623489882E8, 9.623489892E8, 9.623489902E8, 9.623489912E8, 9.623489922E8, 9.623489932E8, 9.623489942E8, 9.623489952E8, 9.623489962E8, 9.623489972E8, 9.623489982E8, 9.623489992E8, 9.623490002E8, 9.623490012E8, 9.623490022E8, 9.623490032E8, 9.623490042E8, 9.623490052E8, 9.623490062E8, 9.623490072E8, 9.623490082E8, 9.623490092E8, 9.623490102E8, 9.623490112E8, 9.623490117E8, 9.623490127E8, 9.623490137E8, 9.623490147E8, 9.623490157E8, 9.623490167E8, 9.623490177E8, 9.623490187E8, 9.623490197E8, 9.623490207E8, 9.623490218E8, 9.623490228E8, 9.623490238E8, 9.623490248E8, 9.623490258E8, 9.623490268E8, 9.623490278E8, 9.623490288E8, 9.623490298E8, 9.623490308E8, 9.623490318E8, 9.623490328E8, 9.623490338E8, 9.623490348E8, 9.623490358E8, 9.623490368E8, 9.623490378E8, 9.623490388E8, 9.623490398E8, 9.623490408E8, 9.623490418E8, 9.623490428E8, 9.623490438E8, 9.623490448E8, 9.623490458E8, 9.623490468E8, 9.623490478E8, 9.623490488E8, 9.623490498E8, 9.623490508E8, 9.623490518E8, 9.623490528E8, 9.623490538E8, 9.623490548E8, 9.623490558E8, 9.623490568E8, 9.623490578E8, 9.623490588E8, 9.623490598E8, 9.623490608E8, 9.623490618E8, 9.623490628E8, 9.623490638E8, 9.623490648E8, 9.623490658E8, 9.623490668E8, 9.623490678E8, 9.623490688E8, 9.623490698E8, 9.623490708E8, 9.623490718E8, 9.623490723E8, 9.623490733E8, 9.623490743E8, 9.623490753E8, 9.623490763E8, 9.623490773E8, 9.623490783E8, 9.623490793E8, 9.623490803E8, 9.623490813E8, 9.623490823E8, 9.623490833E8, 9.623490843E8, 9.623490853E8, 9.623490863E8, 9.623490873E8, 9.623490883E8, 9.623490893E8, 9.623490903E8, 9.623490913E8, 9.623490923E8, 9.623490933E8, 9.623490943E8, 9.623490953E8, 9.623490963E8, 9.623490973E8, 9.623490983E8, 9.623490993E8, 9.623491003E8, 9.623491013E8, 9.623491023E8, 9.623491033E8, 9.623491043E8, 9.623491053E8, 9.623491063E8, 9.623491073E8, 9.623491083E8, 9.623491093E8, 9.623491103E8, 9.623491113E8, 9.623491123E8, 9.623491133E8, 9.623491138E8, 9.623491148E8, 9.623491158E8, 9.623491168E8, 9.623491178E8, 9.623491188E8, 9.623491198E8, 9.623491208E8, 9.623491218E8, 9.623491228E8, 9.623491239E8, 9.623491249E8, 9.623491259E8, 9.623491269E8, 9.623491279E8, 9.623491289E8, 9.623491299E8, 9.623491309E8, 9.623491319E8, 9.623491329E8, 9.623491339E8, 9.623491349E8, 9.623491359E8, 9.623491369E8, 9.623491379E8, 9.623491389E8, 9.623491399E8, 9.623491409E8, 9.623491419E8, 9.623491429E8, 9.623491439E8, 9.623491449E8, 9.623491459E8, 9.623491469E8, 9.623491479E8, 9.623491489E8, 9.623491499E8, 9.623491509E8, 9.623491519E8, 9.623491529E8, 9.623491539E8, 9.623491549E8, 9.623491559E8, 9.623491569E8, 9.623491579E8, 9.623491589E8, 9.623491599E8, 9.623491609E8, 9.623491619E8, 9.623491629E8, 9.623491639E8, 9.623491649E8, 9.623491659E8, 9.623491669E8, 9.623491679E8, 9.623491689E8, 9.623491699E8, 9.623491709E8, 9.623491719E8, 9.623491729E8, 9.623491739E8, 9.623491749E8, 9.623491759E8, 9.623491769E8, 9.623491779E8, 9.623491789E8, 9.623491799E8, 9.623491809E8, 9.623491819E8, 9.623491829E8, 9.623491839E8, 9.623491849E8, 9.623491859E8, 9.623491869E8, 9.623491879E8, 9.623491889E8, 9.623491899E8, 9.623491909E8, 9.623491919E8, 9.623491929E8, 9.623491939E8, 9.623491949E8, 9.623491959E8, 9.623491969E8, 9.623491979E8, 9.623491989E8, 9.623491999E8, 9.623492009E8, 9.623492019E8, 9.623492029E8, 9.623492039E8, 9.623492049E8, 9.623492059E8, 9.623492069E8, 9.623492079E8, 9.623492089E8, 9.623492099E8, 9.623492109E8, 9.623492119E8, 9.623492129E8, 9.623492139E8, 9.623492149E8, 9.623492154E8, 9.623492164E8, 9.623492174E8, 9.623492184E8, 9.623492194E8, 9.623492204E8, 9.623492214E8, 9.623492224E8, 9.623492234E8, 9.623492244E8, 9.623492255E8, 9.623492265E8, 9.623492275E8, 9.623492285E8, 9.623492295E8, 9.623492305E8, 9.623492315E8, 9.623492325E8, 9.623492335E8, 9.623492345E8, 9.623492355E8, 9.623492365E8, 9.623492375E8, 9.623492385E8, 9.623492395E8, 9.623492405E8, 9.623492415E8, 9.623492425E8, 9.623492435E8, 9.623492445E8, 9.623492455E8, 9.623492465E8, 9.623492475E8, 9.623492485E8, 9.623492495E8, 9.623492505E8, 9.623492515E8, 9.623492525E8, 9.623492535E8, 9.623492545E8, 9.623492555E8, 9.623492565E8, 9.623492575E8, 9.623492585E8, 9.623492595E8, 9.623492605E8, 9.623492615E8, 9.623492625E8, 9.623492635E8, 9.623492645E8, 9.623492655E8, 9.623492665E8, 9.623492675E8, 9.623492685E8, 9.623492695E8, 9.623492705E8, 9.623492715E8, 9.623492725E8, 9.623492735E8, 9.623492745E8, 9.623492755E8, 9.623492765E8, 9.623492775E8, 9.623492785E8, 9.623492795E8, 9.623492805E8, 9.623492815E8, 9.623492825E8, 9.623492835E8, 9.623492845E8, 9.623492855E8, 9.623492865E8, 9.623492875E8, 9.623492885E8, 9.623492895E8, 9.623492905E8, 9.623492915E8, 9.623492925E8, 9.623492935E8, 9.623492945E8, 9.623492955E8, 9.623492965E8, 9.62349297E8, 9.62349298E8, 9.62349299E8, 9.623493E8, 9.62349301E8, 9.62349302E8, 9.62349303E8, 9.62349304E8, 9.62349305E8, 9.62349306E8, 9.62349307E8, 9.62349308E8, 9.62349309E8, 9.6234931E8, 9.62349311E8, 9.62349312E8, 9.62349313E8, 9.62349314E8, 9.62349315E8, 9.62349316E8, 9.62349317E8, 9.62349318E8, 9.62349319E8, 9.6234932E8, 9.62349321E8, 9.62349322E8, 9.62349323E8, 9.62349324E8, 9.62349325E8, 9.62349326E8, 9.62349327E8, 9.62349328E8, 9.62349329E8, 9.6234933E8, 9.62349331E8, 9.62349332E8, 9.62349333E8, 9.62349334E8, 9.62349335E8, 9.62349336E8, 9.62349337E8, 9.623493381E8, 9.623493391E8, 9.623493401E8, 9.623493411E8, 9.623493421E8, 9.623493431E8, 9.623493441E8, 9.623493451E8, 9.623493461E8, 9.623493471E8, 9.623493481E8, 9.623493491E8, 9.623493501E8, 9.623493511E8, 9.623493521E8, 9.623493531E8, 9.623493541E8, 9.623493551E8, 9.623493561E8, 9.623493571E8, 9.623493581E8, 9.623493591E8, 9.623493601E8, 9.623493611E8, 9.623493621E8, 9.623493631E8, 9.623493641E8, 9.623493651E8, 9.623493661E8, 9.623493671E8, 9.623493681E8, 9.623493691E8, 9.623493701E8, 9.623493711E8, 9.623493721E8, 9.623493731E8, 9.623493741E8, 9.623493751E8, 9.623493761E8, 9.623493771E8, 9.623493781E8, 9.623493791E8, 9.623493801E8, 9.623493811E8, 9.623493821E8, 9.623493831E8, 9.623493841E8, 9.623493851E8, 9.623493861E8, 9.623493871E8, 9.623493881E8, 9.623493891E8, 9.623493901E8, 9.623493911E8, 9.623493921E8, 9.623493931E8, 9.623493941E8, 9.623493951E8, 9.623493961E8, 9.623493971E8, 9.623493981E8, 9.623493991E8, 9.623494001E8, 9.623494011E8, 9.623494021E8, 9.623494031E8, 9.623494041E8, 9.623494051E8, 9.623494061E8, 9.623494071E8, 9.623494081E8, 9.623494091E8, 9.623494101E8, 9.623494111E8, 9.623494121E8, 9.623494131E8, 9.623494141E8, 9.623494151E8, 9.623494161E8, 9.623494171E8, 9.623494181E8, 9.623494191E8, 9.623494201E8, 9.623494211E8, 9.623494221E8, 9.623494231E8, 9.623494241E8, 9.623494251E8, 9.623494261E8, 9.623494271E8, 9.623494281E8, 9.623494291E8, 9.623494301E8, 9.623494311E8, 9.623494321E8, 9.623494331E8, 9.623494341E8, 9.623494351E8, 9.623494361E8, 9.623494371E8, 9.623494381E8, 9.623494391E8, 9.623494402E8, 9.623494412E8, 9.623494422E8, 9.623494432E8, 9.623494442E8, 9.623494452E8, 9.623494462E8, 9.623494472E8, 9.623494482E8, 9.623494492E8, 9.623494502E8, 9.623494512E8, 9.623494522E8, 9.623494532E8, 9.623494542E8, 9.623494552E8, 9.623494562E8, 9.623494572E8, 9.623494582E8, 9.623494592E8, 9.623494602E8, 9.623494612E8, 9.623494622E8, 9.623494632E8, 9.623494642E8, 9.623494652E8, 9.623494662E8, 9.623494672E8, 9.623494682E8, 9.623494692E8, 9.623494702E8, 9.623494712E8, 9.623494722E8, 9.623494732E8, 9.623494742E8, 9.623494752E8, 9.623494762E8, 9.623494772E8, 9.623494782E8, 9.623494792E8, 9.623494802E8, 9.623494812E8, 9.623494822E8, 9.623494832E8, 9.623494842E8, 9.623494852E8, 9.623494862E8, 9.623494872E8, 9.623494882E8, 9.623494892E8, 9.623494902E8, 9.623494912E8, 9.623494922E8, 9.623494932E8, 9.623494942E8, 9.623494952E8, 9.623494962E8, 9.623494972E8, 9.623494982E8, 9.623494992E8, 9.623495002E8, 9.623495012E8, 9.623495022E8, 9.623495032E8, 9.623495042E8, 9.623495052E8, 9.623495062E8, 9.623495072E8, 9.623495082E8, 9.623495092E8, 9.623495102E8, 9.623495112E8, 9.623495122E8, 9.623495127E8, 9.623495137E8, 9.623495147E8, 9.623495157E8, 9.623495167E8, 9.623495177E8, 9.623495187E8, 9.623495197E8, 9.623495207E8, 9.623495217E8, 9.623495222E8, 9.623495232E8, 9.623495242E8, 9.623495252E8, 9.623495262E8, 9.623495272E8, 9.623495282E8, 9.623495292E8, 9.623495302E8, 9.623495312E8, 9.623495323E8, 9.623495333E8, 9.623495343E8, 9.623495353E8, 9.623495363E8, 9.623495373E8, 9.623495383E8, 9.623495393E8, 9.623495403E8, 9.623495413E8, 9.623495423E8, 9.623495433E8, 9.623495443E8, 9.623495453E8, 9.623495463E8, 9.623495473E8, 9.623495483E8, 9.623495493E8, 9.623495503E8, 9.623495513E8, 9.623495518E8, 9.623495528E8, 9.623495538E8, 9.623495548E8, 9.623495558E8, 9.623495568E8, 9.623495578E8, 9.623495588E8, 9.623495598E8, 9.623495608E8, 9.623495618E8, 9.623495623E8, 9.623495633E8, 9.623495643E8, 9.623495653E8, 9.623495663E8, 9.623495673E8, 9.623495683E8, 9.623495693E8, 9.623495703E8, 9.623495713E8, 9.623495723E8, 9.623495728E8, 9.623495738E8, 9.623495748E8, 9.623495758E8, 9.623495768E8, 9.623495778E8, 9.623495788E8, 9.623495798E8, 9.623495808E8, 9.623495818E8, 9.623495828E8, 9.623495838E8, 9.623495848E8, 9.623495858E8, 9.623495868E8, 9.623495878E8, 9.623495888E8, 9.623495898E8, 9.623495908E8, 9.623495918E8, 9.623495928E8, 9.623495938E8, 9.623495948E8, 9.623495958E8, 9.623495968E8, 9.623495978E8, 9.623495988E8, 9.623495998E8, 9.623496008E8, 9.623496018E8, 9.623496028E8, 9.623496038E8, 9.623496048E8, 9.623496058E8, 9.623496068E8, 9.623496078E8, 9.623496088E8, 9.623496098E8, 9.623496108E8, 9.623496118E8, 9.623496128E8, 9.623496138E8, 9.623496143E8, 9.623496153E8, 9.623496163E8, 9.623496173E8, 9.623496183E8, 9.623496193E8, 9.623496203E8, 9.623496213E8, 9.623496223E8, 9.623496233E8, 9.623496238E8, 9.623496248E8, 9.623496258E8, 9.623496268E8, 9.623496278E8, 9.623496288E8, 9.623496298E8, 9.623496308E8, 9.623496318E8, 9.623496328E8, 9.623496338E8, 9.623496343E8, 9.623496353E8, 9.623496363E8, 9.623496373E8, 9.623496383E8, 9.623496393E8, 9.623496403E8, 9.623496413E8, 9.623496423E8, 9.623496428E8, 9.623496438E8, 9.623496444E8, 9.623496454E8, 9.623496464E8, 9.623496474E8, 9.623496484E8, 9.623496494E8, 9.623496504E8, 9.623496514E8, 9.623496524E8, 9.623496534E8, 9.623496544E8, 9.623496554E8, 9.623496564E8, 9.623496574E8, 9.623496584E8, 9.623496594E8, 9.623496604E8, 9.623496614E8, 9.623496624E8, 9.623496634E8, 9.623496644E8, 9.623496654E8, 9.623496664E8, 9.623496674E8, 9.623496684E8, 9.623496694E8, 9.623496704E8, 9.623496714E8, 9.623496724E8, 9.623496734E8, 9.623496744E8, 9.623496749E8, 9.623496759E8, 9.623496769E8, 9.623496779E8, 9.623496789E8, 9.623496799E8, 9.623496809E8, 9.623496819E8, 9.623496829E8, 9.623496839E8, 9.623496849E8, 9.623496859E8, 9.623496869E8, 9.623496879E8, 9.623496889E8, 9.623496899E8, 9.623496909E8, 9.623496919E8, 9.623496929E8, 9.623496939E8, 9.623496949E8, 9.623496959E8, 9.623496969E8, 9.623496979E8, 9.623496989E8, 9.623496999E8, 9.623497009E8, 9.623497019E8, 9.623497029E8, 9.623497039E8, 9.623497049E8, 9.623497059E8, 9.623497069E8, 9.623497079E8, 9.623497089E8, 9.623497099E8, 9.623497109E8, 9.623497119E8, 9.623497129E8, 9.623497139E8, 9.623497149E8, 9.623497154E8, 9.623497164E8, 9.623497174E8, 9.623497184E8, 9.623497194E8, 9.623497204E8, 9.623497214E8, 9.623497224E8, 9.623497234E8, 9.623497244E8, 9.623497254E8, 9.623497264E8, 9.623497274E8, 9.623497284E8, 9.623497294E8, 9.623497304E8, 9.623497314E8, 9.623497324E8, 9.623497334E8, 9.623497344E8, 9.623497355E8, 9.623497365E8, 9.623497375E8, 9.623497385E8, 9.623497395E8, 9.623497405E8, 9.623497415E8, 9.623497425E8, 9.623497435E8, 9.623497445E8, 9.623497455E8, 9.623497465E8, 9.623497475E8, 9.623497485E8, 9.623497495E8, 9.623497505E8, 9.623497515E8, 9.623497525E8, 9.623497535E8, 9.623497545E8, 9.623497555E8, 9.623497565E8, 9.62349757E8, 9.62349758E8, 9.62349759E8, 9.6234976E8, 9.62349761E8, 9.62349762E8, 9.62349763E8, 9.62349764E8, 9.62349765E8, 9.62349766E8, 9.62349767E8, 9.62349768E8, 9.62349769E8, 9.6234977E8, 9.62349771E8, 9.62349772E8, 9.62349773E8, 9.62349774E8, 9.62349775E8, 9.62349776E8, 9.62349777E8, 9.62349778E8, 9.62349779E8, 9.6234978E8, 9.62349781E8, 9.62349782E8, 9.62349783E8, 9.62349784E8, 9.62349785E8, 9.62349786E8, 9.62349787E8, 9.62349788E8, 9.62349789E8, 9.6234979E8, 9.62349791E8, 9.62349792E8, 9.62349793E8, 9.62349794E8, 9.62349795E8, 9.62349796E8, 9.62349797E8, 9.62349798E8, 9.623497985E8, 9.623497995E8, 9.623498005E8, 9.623498015E8, 9.623498025E8, 9.623498035E8, 9.623498045E8, 9.623498055E8, 9.623498065E8, 9.623498075E8, 9.623498085E8, 9.623498095E8, 9.623498105E8, 9.623498115E8, 9.623498125E8, 9.623498135E8, 9.623498145E8, 9.623498155E8, 9.623498165E8, 9.623498175E8, 9.623498185E8, 9.623498195E8, 9.623498205E8, 9.623498215E8, 9.623498225E8, 9.623498235E8, 9.623498245E8, 9.623498255E8, 9.623498265E8, 9.623498275E8, 9.623498285E8, 9.623498295E8, 9.623498305E8, 9.623498315E8, 9.623498325E8, 9.623498335E8, 9.623498345E8, 9.623498355E8, 9.623498365E8, 9.623498376E8, 9.623498386E8, 9.623498396E8, 9.623498406E8, 9.623498416E8, 9.623498426E8, 9.623498436E8, 9.623498446E8, 9.623498456E8, 9.623498466E8, 9.623498476E8, 9.623498486E8, 9.623498491E8, 9.623498501E8, 9.623498511E8, 9.623498521E8, 9.623498531E8, 9.623498541E8, 9.623498551E8, 9.623498561E8, 9.623498571E8, 9.623498581E8, 9.623498591E8, 9.623498601E8, 9.623498611E8, 9.623498621E8, 9.623498631E8, 9.623498641E8, 9.623498651E8, 9.623498661E8, 9.623498671E8, 9.623498681E8, 9.623498691E8, 9.623498701E8, 9.623498711E8, 9.623498721E8, 9.623498731E8, 9.623498741E8, 9.623498751E8, 9.623498761E8, 9.623498771E8, 9.623498781E8, 9.623498791E8, 9.623498801E8, 9.623498811E8, 9.623498821E8, 9.623498831E8, 9.623498841E8, 9.623498851E8, 9.623498861E8, 9.623498871E8, 9.623498881E8, 9.623498891E8, 9.623498901E8, 9.623498911E8, 9.623498921E8, 9.623498931E8, 9.623498941E8, 9.623498951E8, 9.623498961E8, 9.623498971E8, 9.623498981E8, 9.623498991E8, 9.623498996E8, 9.623499006E8, 9.623499016E8, 9.623499026E8, 9.623499036E8, 9.623499046E8, 9.623499056E8, 9.623499066E8, 9.623499076E8, 9.623499086E8, 9.623499096E8, 9.623499106E8, 9.623499116E8, 9.623499126E8, 9.623499136E8, 9.623499146E8, 9.623499156E8, 9.623499166E8, 9.623499176E8, 9.623499186E8, 9.623499196E8, 9.623499201E8, 9.623499211E8, 9.623499221E8, 9.623499231E8, 9.623499241E8, 9.623499251E8, 9.623499261E8, 9.623499271E8, 9.623499281E8, 9.623499291E8, 9.623499301E8, 9.623499311E8, 9.623499321E8, 9.623499331E8, 9.623499341E8, 9.623499351E8, 9.623499361E8, 9.623499371E8, 9.623499381E8, 9.623499391E8, 9.623499401E8, 9.623499411E8, 9.623499421E8, 9.623499431E8, 9.623499441E8, 9.623499451E8, 9.623499461E8, 9.623499471E8, 9.623499481E8, 9.623499491E8, 9.623499502E8, 9.623499512E8, 9.623499522E8, 9.623499532E8, 9.623499542E8, 9.623499552E8, 9.623499562E8, 9.623499572E8, 9.623499582E8, 9.623499592E8, 9.623499602E8, 9.623499612E8, 9.623499622E8, 9.623499632E8, 9.623499642E8, 9.623499652E8, 9.623499662E8, 9.623499672E8, 9.623499682E8, 9.623499692E8, 9.623499702E8, 9.623499712E8, 9.623499717E8, 9.623499727E8, 9.623499737E8, 9.623499747E8, 9.623499757E8, 9.623499767E8, 9.623499777E8, 9.623499787E8, 9.623499797E8, 9.623499807E8, 9.623499817E8, 9.623499827E8, 9.623499837E8, 9.623499847E8, 9.623499857E8, 9.623499867E8, 9.623499877E8, 9.623499887E8, 9.623499897E8, 9.623499907E8, 9.623499917E8, 9.623499927E8, 9.623499937E8, 9.623499947E8, 9.623499957E8, 9.623499967E8, 9.623499977E8, 9.623499987E8, 9.623499997E8, 9.623500007E8, 9.623500017E8, 9.623500027E8, 9.623500032E8, 9.623500042E8, 9.623500052E8, 9.623500062E8, 9.623500072E8, 9.623500082E8, 9.623500092E8, 9.623500102E8, 9.623500112E8, 9.623500117E8, 9.623500127E8, 9.623500137E8, 9.623500147E8, 9.623500157E8, 9.623500167E8, 9.623500177E8, 9.623500187E8, 9.623500197E8, 9.623500207E8, 9.623500217E8, 9.623500222E8, 9.623500232E8, 9.623500242E8, 9.623500252E8, 9.623500262E8, 9.623500272E8, 9.623500282E8, 9.623500292E8, 9.623500302E8, 9.623500312E8, 9.623500322E8, 9.623500327E8, 9.623500337E8, 9.623500347E8, 9.623500357E8, 9.623500367E8, 9.623500377E8, 9.623500387E8, 9.623500397E8, 9.623500407E8, 9.623500418E8, 9.623500428E8, 9.623500438E8, 9.623500448E8, 9.623500458E8, 9.623500468E8, 9.623500478E8, 9.623500488E8, 9.623500498E8, 9.623500508E8, 9.623500518E8, 9.623500528E8, 9.623500533E8, 9.623500543E8, 9.623500553E8, 9.623500563E8, 9.623500573E8, 9.623500583E8, 9.623500593E8, 9.623500603E8, 9.623500613E8, 9.623500623E8, 9.623500633E8, 9.623500638E8, 9.623500648E8, 9.623500658E8, 9.623500668E8, 9.623500678E8, 9.623500688E8, 9.623500698E8, 9.623500708E8, 9.623500718E8, 9.623500728E8, 9.623500738E8, 9.623500743E8, 9.623500753E8, 9.623500763E8, 9.623500773E8, 9.623500783E8, 9.623500793E8, 9.623500803E8, 9.623500813E8, 9.623500823E8, 9.623500833E8, 9.623500838E8, 9.623500848E8, 9.623500858E8, 9.623500868E8, 9.623500878E8, 9.623500888E8, 9.623500898E8, 9.623500908E8, 9.623500918E8, 9.623500928E8, 9.623500938E8, 9.623500948E8, 9.623500958E8, 9.623500968E8, 9.623500978E8, 9.623500988E8, 9.623500998E8, 9.623501008E8, 9.623501018E8, 9.623501028E8, 9.623501038E8, 9.623501043E8, 9.623501053E8, 9.623501063E8, 9.623501073E8, 9.623501083E8, 9.623501093E8, 9.623501103E8, 9.623501113E8, 9.623501123E8, 9.623501133E8, 9.623501143E8, 9.623501153E8, 9.623501163E8, 9.623501173E8, 9.623501183E8, 9.623501193E8, 9.623501203E8, 9.623501213E8, 9.623501223E8, 9.623501233E8, 9.623501243E8, 9.623501253E8, 9.623501263E8, 9.623501273E8, 9.623501283E8, 9.623501293E8, 9.623501303E8, 9.623501313E8, 9.623501323E8, 9.623501333E8, 9.623501343E8, 9.623501348E8, 9.623501358E8, 9.623501368E8, 9.623501378E8, 9.623501388E8, 9.623501398E8, 9.623501408E8, 9.623501418E8, 9.623501428E8, 9.623501438E8, 9.623501443E8, 9.623501453E8, 9.623501463E8, 9.623501473E8, 9.623501483E8, 9.623501493E8, 9.623501503E8, 9.623501513E8, 9.623501523E8, 9.623501533E8, 9.623501544E8, 9.623501554E8, 9.623501564E8, 9.623501574E8, 9.623501584E8, 9.623501594E8, 9.623501604E8, 9.623501614E8, 9.623501624E8, 9.623501634E8, 9.623501644E8, 9.623501649E8, 9.623501659E8, 9.623501669E8, 9.623501679E8, 9.623501689E8, 9.623501699E8, 9.623501709E8, 9.623501719E8, 9.623501729E8, 9.623501739E8, 9.623501749E8, 9.623501754E8, 9.623501764E8, 9.623501774E8, 9.623501784E8, 9.623501794E8, 9.623501804E8, 9.623501814E8, 9.623501824E8, 9.623501834E8, 9.623501844E8, 9.623501854E8, 9.623501859E8, 9.623501869E8, 9.623501879E8, 9.623501889E8, 9.623501899E8, 9.623501909E8, 9.623501919E8, 9.623501929E8, 9.623501939E8, 9.623501949E8, 9.623501959E8, 9.623501964E8, 9.623501974E8, 9.623501984E8, 9.623501994E8, 9.623502004E8, 9.623502014E8, 9.623502024E8, 9.623502034E8, 9.623502044E8, 9.623502054E8, 9.623502064E8, 9.623502069E8, 9.623502079E8, 9.623502089E8, 9.623502099E8, 9.623502109E8, 9.623502119E8, 9.623502129E8, 9.623502139E8, 9.623502149E8, 9.623502159E8, 9.623502169E8, 9.623502179E8, 9.623502189E8, 9.623502199E8, 9.623502209E8, 9.623502219E8, 9.623502229E8, 9.623502239E8, 9.623502249E8, 9.623502259E8, 9.623502269E8, 9.623502279E8, 9.623502289E8, 9.623502299E8, 9.623502309E8, 9.623502319E8, 9.623502329E8, 9.623502339E8, 9.623502349E8, 9.623502359E8, 9.623502369E8, 9.623502374E8, 9.623502384E8, 9.623502394E8, 9.623502404E8, 9.623502414E8, 9.623502424E8, 9.623502434E8, 9.623502444E8, 9.623502454E8, 9.623502465E8, 9.623502475E8, 9.623502485E8, 9.623502495E8, 9.623502505E8, 9.623502515E8, 9.623502525E8, 9.623502535E8, 9.623502545E8, 9.623502555E8, 9.623502565E8, 9.62350257E8, 9.62350258E8, 9.62350259E8, 9.6235026E8, 9.62350261E8, 9.62350262E8, 9.62350263E8, 9.62350264E8, 9.62350265E8, 9.62350266E8, 9.62350267E8, 9.62350268E8, 9.62350269E8, 9.6235027E8, 9.62350271E8, 9.62350272E8, 9.62350273E8, 9.62350274E8, 9.62350275E8, 9.62350276E8, 9.62350277E8, 9.623502775E8, 9.623502785E8, 9.623502795E8, 9.623502805E8, 9.623502815E8, 9.623502825E8, 9.623502835E8, 9.623502845E8, 9.623502855E8, 9.623502865E8, 9.62350287E8, 9.62350288E8, 9.62350289E8, 9.6235029E8, 9.62350291E8, 9.62350292E8, 9.62350293E8, 9.62350294E8, 9.62350295E8, 9.62350296E8, 9.62350297E8, 9.62350298E8, 9.623502985E8, 9.623502995E8, 9.623503005E8, 9.623503015E8, 9.623503025E8, 9.623503035E8, 9.623503045E8, 9.623503055E8, 9.623503065E8, 9.623503075E8, 9.623503085E8, 9.623503095E8, 9.623503105E8, 9.623503115E8, 9.623503125E8, 9.623503135E8, 9.623503145E8, 9.623503155E8, 9.623503165E8, 9.623503175E8, 9.62350318E8, 9.62350319E8, 9.6235032E8, 9.62350321E8, 9.62350322E8, 9.62350323E8, 9.62350324E8, 9.62350325E8, 9.62350326E8, 9.62350327E8, 9.62350328E8, 9.62350329E8, 9.623503295E8, 9.623503305E8, 9.623503315E8, 9.623503325E8, 9.623503335E8, 9.623503345E8, 9.623503355E8, 9.623503365E8, 9.623503375E8, 9.623503385E8, 9.623503395E8, 9.623503405E8, 9.623503415E8, 9.623503425E8, 9.623503435E8, 9.623503445E8, 9.623503455E8, 9.623503465E8, 9.623503475E8, 9.623503485E8, 9.623503491E8, 9.623503501E8, 9.623503511E8, 9.623503521E8, 9.623503531E8, 9.623503541E8, 9.623503551E8, 9.623503561E8, 9.623503571E8, 9.623503581E8, 9.623503586E8, 9.623503596E8, 9.623503606E8, 9.623503616E8, 9.623503626E8, 9.623503636E8, 9.623503646E8, 9.623503656E8, 9.623503666E8, 9.623503676E8, 9.623503686E8, 9.623503696E8, 9.623503706E8, 9.623503716E8, 9.623503726E8, 9.623503736E8, 9.623503746E8, 9.623503756E8, 9.623503766E8, 9.623503776E8, 9.623503786E8, 9.623503791E8, 9.623503801E8, 9.623503811E8, 9.623503821E8, 9.623503831E8, 9.623503841E8, 9.623503851E8, 9.623503861E8, 9.623503871E8, 9.623503881E8, 9.623503891E8, 9.623503901E8, 9.623503911E8, 9.623503921E8, 9.623503931E8, 9.623503941E8, 9.623503951E8, 9.623503961E8, 9.623503971E8, 9.623503981E8, 9.623503991E8, 9.623504001E8, 9.623504011E8, 9.623504021E8, 9.623504031E8, 9.623504041E8, 9.623504051E8, 9.623504061E8, 9.623504071E8, 9.623504081E8, 9.623504091E8, 9.623504101E8, 9.623504111E8, 9.623504116E8, 9.623504126E8, 9.623504136E8, 9.623504146E8, 9.623504156E8}
pres =
  {898.5, -999.0, -999.0, -999.0, -999.0, -999.0, 898.3279, 897.96155, 897.58875, 897.2087, 896.8203, 896.42255, 896.0142, 895.59454, 895.1633, 894.7208, 894.26715, 893.80273, 893.3284, 892.8454, 892.35474, 891.85754, 891.35474, 890.8473, 890.3361, 889.8222, 889.3066, 888.7903, 888.2745, 887.7602, 887.2484, 886.74005, 886.2361, 885.7374, 885.24506, 884.75977, 884.28253, 883.8142, 883.35547, 882.907, 882.4694, 882.0432, 881.6285, 881.225, 880.8326, 880.45105, 880.08, 879.719, 879.3677, 879.0256, 878.6923, 878.3677, 878.05133, 877.74286, 877.4416, 877.14636, 876.8564, 876.5706, 876.28845, 876.0094, 875.7053, 875.43115, 875.1594, 874.89087, 874.6259, 874.3652, 874.1087, 873.85645, 873.6085, 873.36487, 873.1254, 872.8904, 872.65967, 872.4335, 872.2129, 871.9993, 871.79395, 871.59814, 871.41315, 871.24023, 871.08075, 870.9358, 870.8061, 870.69226, 870.59503, 870.5146, 870.4503, 870.401, 870.3656, 870.3429, 870.33075, 870.32684, -999.0, -999.0, -999.0, -999.0, -999.0, 870.3065, 870.26624, 870.20416, 870.1162, 869.9986, 869.8493, 869.6669, 869.4498, 869.197, 868.909, 868.58673, 868.2312, 867.8436, 867.4262, 866.98145, 866.5117, 866.0196, 865.5077, 864.9786, 864.4349, 863.8794, 863.31506, 862.74493, 862.17206, 861.5993, 861.02924, 860.4639, 859.9057, 859.3566, 858.818, 858.2907, 857.77594, 857.2746, 856.78766, 856.3159, 855.8603, 855.4215, 854.99963, 854.5946, 854.2063, 853.83453, 853.47864, 853.13794, 852.81165, 852.4991, 852.1991, 851.9106, 851.6325, 851.36346, 851.1017, 850.84503, 850.59143, 850.33887, 850.08563, 849.83014, 849.57086, 849.3062, 849.0355, 848.7583, 848.474, 848.18225, 847.88354, 847.5477, 847.23676, 846.92114, 846.60223, 846.2815, 845.9603, 845.6401, 845.32117, 845.004, 844.68896, 844.3762, 844.06537, 843.75586, 843.4471, 843.13855, 842.82947, 842.5191, 842.20654, 841.8912, 841.5723, 841.24945, 840.9221, 840.5898, 840.2518, 839.90753, 839.5565, 839.19806, 838.8315, 838.4559, 838.07043, 837.6745, 837.26776, 836.85016, 836.4214, 835.98175, 835.5324, 835.075, 834.6112, 834.1427, 833.67163, 833.2002, 832.7306, 832.2649, 831.8046, 831.3511, 830.90564, 830.4696, 830.04376, 829.629, 829.2261, 828.8357, 828.4582, 828.09375, 827.74255, 827.4046, 827.0792, 826.7653, 826.462, 826.168, 825.88196, 825.60205, 825.32654, 825.0538, 824.78253, 824.51166, 824.24, 823.9666, 823.6909, 823.4126, 823.13135, 822.8469, 822.55927, 822.26843, 821.9745, 821.6777, 821.3784, 821.07745, 820.7754, 820.4729, 820.1709, 819.8702, 819.57153, 819.276, 818.9845, 818.6981, 818.41797, 818.14496, 817.8796, 817.62213, 817.3728, 817.13184, 816.89886, 816.67334, 816.4548, 816.2426, 816.036, 815.83417, 815.63617, 815.4411, 815.24817, 815.05646, 814.8651, 814.6733, 814.4804, 814.26654, 814.0701, 813.8716, 813.67114, 813.46936, 813.2667, 813.06384, 812.86176, 812.6617, 812.4648, 812.27234, 812.08527, 811.9044, 811.7308, 811.5651, 811.4082, 811.26044, 811.1225, 810.99493, 810.8783, 810.77325, 810.6803, 810.6001, 810.5329, 810.4792, 810.43915, 810.413, 810.4007, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 810.33966, 810.1036, 809.8599, 809.6077, 809.3457, 809.0726, 808.78705, 808.4571, 808.1416, 807.81036, 807.4626, 807.09735, 806.7144, 806.3136, 805.8948, 805.4579, 805.00354, 804.5324, 804.0453, 803.5429, 803.0264, 802.49713, 801.9562, 801.4049, 800.8449, 800.2781, 799.70605, 799.13074, 798.5539, 797.97754, 797.4034, 796.8334, 796.2691, 795.7121, 795.1639, 794.626, 794.0994, 793.5851, 793.08405, 792.597, 792.1239, 791.6645, 791.21844, 790.78546, 790.365, 789.9566, 789.5597, 789.17377, 788.79803, 788.4315, 788.0734, 787.7229, 787.3789, 787.0406, 786.707, 786.37714, 786.0503, 785.7257, 785.40265, 785.0804, 784.75836, 784.43616, 784.1132, 783.7891, 783.46356, 783.1364, 782.80756, 782.47687, 782.14453, 781.8108, 781.47595, 781.1403, 780.8038, 780.46606, 780.1271, 779.78644, 779.4435, 779.0974, 778.7474, 778.39246, 778.0318, 777.6644, 777.2893, 776.90546, 776.51196, 776.10754, 775.6913, 775.26215, 774.8193, 774.36224, 773.8904, 773.4032, 772.9007, 772.3829, 771.8499, 771.302, 770.7398, 770.1641, 769.5759, 768.9154, 768.3035, 767.6816, 767.05023, 766.4103, 765.76263, 765.1083, 764.44806, 763.78296, 763.1143, 762.44324, 761.7711, 761.0991, 760.42847, 759.7603, 759.09576, 758.4359, 757.7813, 757.13226, 756.4891, 755.852, 755.22095, 754.59564, 753.9757, 753.3609, 752.75037, 752.1434, 751.5389, 750.93616, 750.3348, 749.73456, 749.13513, 748.53644, 747.9385, 747.3415, 746.74567, 746.1512, 745.5579, 744.9658, 744.3746, 743.7842, 743.19446, 742.60535, 742.01666, 741.42834, 740.84033, 740.25256, 739.665, 739.0775, 738.49023, 737.9033, 737.3168, 736.7309, 736.1459, 735.5621, 734.98, 734.39984, 733.8219, 733.2464, 732.6735, 732.10345, 731.53595, 730.9705, 730.4068, 729.84424, 729.2823, 728.72, 728.15656, 727.5911, 727.02277, 726.45056, 725.8735, 725.2906, 724.7014, 724.10583, 723.5036, 722.89453, 722.2789, 721.6571, 721.02966, 720.3971, 719.7606, 719.1217, 718.48193, 717.84265, 717.2055, 716.57196, 715.9434, 715.3215, 714.7072, 714.1017, 713.5058, 712.92053, 712.34607, 711.7823, 711.22906, 710.6862, 710.1525, 709.6266, 709.10675, 708.59155, 708.0795, 707.56946, 707.0599, 706.54956, 706.0378, 705.52386, 705.00726, 704.4876, 703.9648, 703.4393, 702.91144, 702.3286, 701.7981, 701.2687, 700.74194, 700.2195, 699.70294, 699.1939, 698.6941, 698.2051, 697.7277, 697.2628, 696.81104, -999.0, -999.0, -999.0, 695.13666, 694.74805, 694.37, 694.0018, 693.64264, 693.2919, 692.94904, 692.61365, 692.2853, 691.96356, 691.64825, 691.33923, 691.03625, 690.7393, 690.44836, 690.1635, 689.8849, 689.6125, 689.3465, 689.0868, 688.83356, 688.58673, 688.3461, 688.1113, 687.8822, 687.65826, 687.43884, 687.2231, 687.01013, 686.7992, 686.58923, 686.37933, 686.16846, 685.9557, 685.74, 685.5204, 685.2958, 685.06525, 684.82825, 684.5844, 684.33344, 684.07513, 683.8098, 683.5383, 683.26135, 682.9796, 682.6935, 682.40314, 682.10864, 681.8102, 681.50745, 681.1999, 680.887, 680.56836, 680.2436, 679.9126, 679.57526, 679.2314, 678.8818, 678.5275, 678.16974, 677.8095, 677.448, 677.0865, 676.72626, 676.36847, 676.0139, 675.6631, 675.31647, 674.9747, 674.63776, 674.3059, 673.9791, 673.6575, 673.34094, 673.02954, 672.7232, 672.392, 672.09625, 671.80554, 671.51984, 671.2391, 670.9627, 670.68976, 670.41956, 670.1512, 669.8834, 669.6151, 669.34503, 669.0719, 668.795, 668.5136, 668.22723, 667.9353, 667.63763, 667.3344, 667.02576, 666.7118, 666.39294, 666.0699, 665.74316, 665.4133, 665.0811, 664.7471, 664.4118, 664.07605, 663.73987, 663.4033, 663.06635, 662.7289, 662.3908, 662.0518, 661.7116, 661.37006, 661.027, 660.6823, 660.3361, 659.9882, 659.6384, 659.28613, 658.93097, 658.5724, 658.20984, 657.8427, 657.4703, 657.09204, 656.70825, 656.3196, 655.9267, 655.5303, 655.1312, 654.7304, 654.32874, 653.9272, 653.52563, 653.12396, 652.72174, 652.3186, 651.9141, 651.50757, 651.0983, 650.68585, 650.2697, 649.8499, 649.42615, 648.9983, 648.56665, 648.13153, 647.6934, 647.2526, 646.8099, 646.36615, 645.9223, 645.4792, 645.03754, 644.59796, 644.1611, 643.7276, 643.2979, 642.87244, 642.45154, 642.0356, 641.62494, 641.2201, 640.8214, 640.4292, 640.0436, 639.6645, 639.2919, 638.92554, 638.56537, 638.211, 637.8621, 637.51843, 637.17975, 636.8461, 636.5175, 636.194, 635.8756, 635.5316, 635.2248, 634.9237, 634.62885, 634.3407, 634.0597, 633.78644, 633.5215, 633.26575, 633.0199, 632.7847, 632.5606, 632.34766, 632.1461, 631.956, 631.7771, 631.6088, 631.45074, 631.30225, 631.1626, 631.0309, 630.90625, 630.7878, 630.6745, 630.56555, 630.46, 630.357, 630.2555, 630.15454, 630.0532, 629.95056, 629.846, 629.739, 629.6291, 629.5159, 629.39923, 629.2791, 629.1555, 629.0285, 628.89825, 628.7651, 628.6293, 628.4911, 628.3511, 628.20966, 628.0674, 627.92487, 627.7824, 627.6404, 627.49915, 627.35895, 627.21985, 627.15063, 627.01294, 626.876, 626.73956, 626.6033, 626.46674, 626.3294, 626.1909, 626.0507, 625.90826, 625.763, 625.61444, 625.4622, 625.306, 625.1455, 624.9805, 624.8112, 624.6379, 624.4606, 624.27966, 624.09515, 623.9073, 623.7162, 623.52203, 623.325, 623.1254, 622.9235, 622.7194, 622.51294, 622.304, 622.0924, 621.87775, 621.6595, 621.4369, 621.20917, 620.97565, 620.7353, 620.48737, 620.23083, 619.9649, 619.6888, 619.40186, 619.1034, 618.79285, 618.4702, 618.1356, 617.78906, 617.4309, 617.0623, 616.6845, 616.2598, 615.8669, 615.4689, 615.06726, 614.66345, 614.25885, 613.85486, 613.45276, 613.05383, 612.6593, 612.2701, 611.8869, 611.5107, 611.1421, 610.7813, 610.42865, 610.08435, 609.7484, 609.42065, 609.1007, 608.7882, 608.4828, 608.18384, 607.8907, 607.6028, 607.3194, 607.0398, 606.7633, 606.4891, 606.21643, 605.945, 605.67426, 605.4037, 605.1329, 604.86127, 604.58844, 604.3137, 604.0369, 603.758, 603.4772, 603.19446, 602.9101, 602.6243, 602.3376, 602.0501, 601.7622, 601.4741, 601.1862, 600.8988, 600.61194, 600.3256, 600.03973, 599.7543, 599.4692, 599.1848, 598.9015, 598.61957, 598.3395, 598.06177, 597.7869, 597.5155, 597.24805, 596.9848, 596.72614, 596.47235, 596.22363, 595.9802, 595.74225, 595.5098, 595.28296, 595.06104, 594.84357, 594.63, 594.4197, 594.21155, 594.00476, 593.79834, 593.5913, 593.383, 593.17267, 592.9597, 592.7434, 592.5233, 592.29913, 592.0704, 591.83673, 591.598, 591.3541, 591.1049, 590.8503, 590.59033, 590.325, 590.05444, 589.7787, 589.49817, 589.21326, 588.92444, 588.632, 588.3366, 588.0388, 587.7392, 587.43823, 587.1056, 586.8018, 586.4967, 586.19037, 585.88306, 585.5751, 585.2667, 584.95825, 584.6501, 584.3425, 584.03595, 583.7305, 583.426, 583.1222, 582.8188, 582.51556, 582.21246, 581.9094, 581.60645, 581.3034, 581.0005, 580.6977, 580.395, 580.09265, 579.79065, 579.4891, 579.18805, 578.88763, 578.5877, 578.2882, 577.98895, 577.68976, 577.39044, 577.0905, 576.7898, 576.48785, 576.1845, 575.8797, 575.57324, 575.2651, 574.9553, 574.7999, 574.48834, 574.1758, 573.8623, 573.5479, 573.2326, 572.9164, 572.59924, 572.28143, 571.963, 571.64417, 571.3252, 571.0064, 570.6881, 570.3707, 570.0543, 569.7391, 569.425, 569.1121, 568.80054, 568.49036, 568.1816, 567.8744, 567.56866, 567.2647, 566.96246, 566.66205, 566.3634, 566.0662, 565.77045, 565.4757, 565.18195, 564.889, 564.5967, 564.3048, 564.0133, 563.72186, 563.4304, 563.13873, 562.8466, 562.5538, 562.26, 561.9651, 561.6689, 561.37164, 561.07336, 560.7742, 560.4743, 560.174, 559.87354, 559.5732, 559.2732, 558.97375, 558.67505, 558.37726, 558.08044, 557.78436, 557.4889, 557.1939, 556.89923, 556.6046, 556.3098, 556.0147, 555.7188, 555.42175, 555.1231, 554.8224, 554.51917, 554.2129, 553.90326, 553.58966, 553.27185, 552.9171, 552.5897, 552.2575, 551.9203, 551.57806, 551.23065, 550.87805, 550.52045, 550.1581, 549.7913, 549.4204, 549.04565, 548.6672, 548.2853, 547.90015, 547.51184, 547.1203, 546.72565, 546.32776, 545.92676, 545.5228, 545.3198, 544.91174, 544.5012, 544.0887, 543.6746, 543.2595, 542.844, 542.4286, 542.01404, 541.60095, 541.1899, 540.7813, 540.3756, 539.973, 539.574, 539.1788, 538.7877, 538.4011, 538.0192, 537.6421, 537.2698, 536.90234, 536.5398, 536.18176, 535.8279, 535.47784, 535.1312, 534.78754, 534.44635, 534.10724, 533.7699, 533.4342, 533.1002, 532.76807, 532.43774, 532.10956, 531.7838, 531.4608, 531.14087, 530.8242, 530.511, 530.2015, 529.8958, 529.5939, 529.2955, 529.0004, 528.70844, 528.4188, 528.1308, 527.8437, 527.5567, 527.2695, 526.98175, 526.69305, 526.4032, 526.11194, 525.81934, 525.5252, 525.2295, 524.93243, 524.63416, 524.3349, 524.0349, 523.73444, 523.4337, 523.1332, 522.833, 522.5331, 522.23334, 521.93365, 521.6338, 521.33356, 521.0324, 520.73016, 520.42633, 520.12054, 519.81244, 519.5016, 519.1877, 518.8705, 518.5498, 518.22546, 518.02905, 517.6987, 517.36487, 517.02765, 516.6874, 516.34436, 515.99927, 515.6527, 515.30524, 514.95746, 514.60986, 514.26294, 513.9172, 513.57294, 513.2306, 512.89044, 512.5528, 512.21783, 511.8859, 511.55707, 511.23163, 510.90967, 510.59116, 510.27618, 509.96475, 509.65677, 509.35196, 509.05014, 508.75107, 508.45456, 508.1604, 507.86835, 507.57822, 507.28976, 507.00266, 506.7166, 506.43137, 506.14664, 505.8622, 505.57782, 505.29324, 505.0085, 504.72372, 504.43906, 504.1547, 503.87088, 503.58792, 503.3061, 503.02573, 502.74704, 502.47018, 502.19525, 501.92236, 501.6514, 501.382, 501.11374, 500.84625, 500.57928, 500.3126, 500.046, 499.7793, 499.51236, 499.24515, 498.9776, 498.70963, 498.44128, 498.17264, 497.9038, 497.6349, 497.36603, 497.0976, 496.8298, 496.56302, 496.29736, 496.0329, 495.7697, 495.50784, 495.24728, 494.98795, 494.7298, 494.47275, 494.21655, 494.08865, 493.83307, 493.57742, 493.32138, 493.06464, 492.80698, 492.54816, 492.28796, 492.02618, 491.7626, 491.4704, 491.20245, 490.9321, 490.65906, 490.38312, 490.1041, 489.82175, 489.5359, 489.24634, 488.953, 488.65585, 488.35498, 488.05048, 487.7424, 487.43103, 487.11664, 486.79944, 486.47977, 486.15784, 485.83398, 485.50848, 485.18164, 484.85394, 484.52594, 484.19818, 483.8712, 483.54562, 483.22214, 482.9014, 482.58395, 482.26984, 481.95898, 481.6513, 481.34674, 481.0451, 480.74615, 480.44968, 480.15546, 479.8632, 479.5726, 479.28333, 478.99512, 478.70767, 478.42072, 478.134, 477.8472, 477.56003, 477.27213, 476.98312, 476.6927, 476.40042, 476.25345, 475.95767, 475.659, 475.3571, 475.0515, 474.74194, 474.42795, 474.1095, 473.78696, 473.46057, 473.13065, 472.7975, 472.46118, 472.12195, 471.77994, 471.43524, 471.08792, 470.738, 470.3855, 470.0304, 469.6726, 469.31198, 468.9485, 468.58188, 468.212, 467.83865, 467.46158, 467.08078, 466.69635, 466.30844, 465.9172, 465.52286, 465.1257, 464.72607, 464.32428, 463.92062, 463.5154, 463.10895, 462.7015, 462.29343, 461.88504, 461.47662, 461.27252, 460.8647, 460.45758, 460.0514, 459.64633, 459.24265, 458.8404, 458.43958, 458.04025, 457.64243, 457.2066, 456.81207, 456.4192, 456.02798, 455.63843, 455.25043, 454.86395, 454.4789, 454.09515, 453.71252, 453.3309, 452.95004, 452.56958, 452.18906, 451.80807, 451.42624, 451.0433, 450.65915, 450.27356, 449.8864, 449.4977, 449.10745, 448.7157, 448.32245, 447.92786, 447.53207, 447.1353, 446.73773, 446.33942, 445.94052, 445.54114, 445.14148, 444.74173, 444.3421, 443.9429, 443.5443, 443.1465, 442.74966, 442.3539, 441.95944, 441.56647, 441.1752, 440.78586, 440.39865, 440.01364, 439.63077, 439.2501, 438.87155, 438.49515, 438.1208, 437.7484, 437.378, 437.0094, 436.64255, 436.2773, 435.9136, 435.5513, 435.1902, 434.8301, 434.47098, 434.11276, 433.7555, 433.3992, 433.04398, 432.68982, 432.3368, 431.98492, 431.6343, 431.28485, 430.93658, 430.58945, 430.2435, 429.8991, 429.55682, 429.21716, 428.88058, 428.54733, 428.21762, 427.89163, 427.5695, 427.25137, 426.93732, 426.6274, 426.32175, 426.0203, 425.723, 425.42984, 425.14075, 424.85562, 424.57437, 424.29688, 424.023, 423.88745, 423.61896, 423.35394, 423.09238, 422.8341, 422.57886, 422.32642, 422.07654, 421.82895, 421.5835, 421.31573, 421.07413, 420.834, 420.59506, 420.35703, 420.11954, 419.8824, 419.64523, 419.40784, 419.16992, 418.93127, 418.6917, 418.45105, 418.20917, 417.96588, 417.72107, 417.4746, 417.22635, 416.9764, 416.7252, 416.47308, 416.22043, 415.96765, 415.71512, 415.46317, 415.21222, 414.96255, 414.71445, 414.46808, 414.2237, 413.98157, 413.74197, 413.50513, 413.2713, 413.0406, 412.8127, 412.58746, 412.3647, 412.14413, 411.92563, 411.70895, 411.49393, 411.28043, 411.0685, 410.85815, 410.6494, 410.4422, 410.23642, 410.03183, 409.82837, 409.62582, 409.4241, 409.22308, 409.02264, 408.82266, 408.62296, 408.42343, 408.2239, 408.02423, 407.82425, 407.62372, 407.42245, 407.22012, 407.01636, 406.8107, 406.60272, 406.39197, 406.178, 405.96042, 405.7387, 405.51245, 405.2811, 405.16333, 404.92337, 404.67703, 404.424, 404.16403, 403.89688, 403.62228, 403.34027, 403.05084, 402.75403, 402.4499, 402.13858, 401.82016, 401.49478, 401.1626, 400.8239, 400.4791, 400.12842, 399.77237, 399.41153, 399.0467, 398.67853, 398.30786, 397.93558, 397.56262, 397.19, 396.81873, 396.45004, 396.0853, 395.72586, 395.37302, 395.02762, 394.6904, 394.36203, 394.04312, 393.73355, 393.43292, 393.14084, 392.8569, 392.58044, 392.31082, 392.0212, 391.76355, 391.51074, 391.2623, 391.01776, 390.7767, 390.53867, 390.30316, 390.06976, 389.838, 389.60742, 389.37756, 389.14798, 388.91818, 388.68784, 388.45663, 388.2242, 387.9903, 387.75485, 387.5179, 387.27957, 387.03983, 386.7987, 386.55627, 386.3126, 386.06766, 385.8216, 385.57443, 385.3263, 385.07724, 384.8272, 384.57614, 384.32397, 384.07068, 383.81638, 383.5612, 383.30533, 383.04895, 382.79193, 382.53418, 382.2756, 382.01605, 381.75543, 381.4937, 381.23077, 380.96658, 380.70117, 380.4345, 380.16672, 379.89777, 379.62775, 379.35678, 379.08493, 378.81232, 378.5391, 378.26553, 377.99185, 377.71823, 377.4447, 377.17133, 376.898, 376.62476, 376.3515, 376.07806, 375.80438, 375.53027, 375.25574, 374.9808, 374.7054, 374.4296, 374.15332, 373.8766, 373.59937, 373.32166, 373.04312, 372.7635, 372.4824, 372.1995, 371.91434, 371.6265, 371.3355, 371.041, 370.74268, 370.44052, 370.13443, 369.82425, 369.51007, 369.1919, 368.86978, 368.54385, 368.21432, 367.8816, 367.546, 367.2079, 366.86777, 366.52618, 366.18365, 365.84076, 365.49792, 365.15567, 364.81442, 364.47464, 364.10306, 363.7676, 363.4348, 363.105, 362.7786, 362.45593, 362.13736, 361.82333, 361.51425, 361.2106, 360.9128, 360.6214, 360.3368, 360.05957, 359.79013, 359.52902, 359.27655, 359.03302, 358.79868, 358.57376, 358.35837, 358.15234, 357.9557, 357.7683, 357.5899, 357.42014, 357.25873, 357.1053, 356.9592, 356.81973, 356.6862, 356.55786, 356.43378, 356.31287, 356.19412, 356.0765, 355.95908, 355.84094, 355.72116, 355.5989, 355.47385, 355.34583, 355.21478, 355.08054, 354.94315, 354.80276, 354.65942, 354.51328, 354.36444, 354.21304, 354.05927, 353.90326, 353.74524, 353.58548, 353.42426, 353.26178, 353.09836, 352.93427, 352.76974, 352.6051, 352.44043, 352.27588, 352.11157, 351.94757, 351.78384, 351.62027, 351.45673, 351.29306, 351.1292, 350.96503, 350.80038, 350.63516, 350.46924, 350.38596, 350.21866, 350.0503, 349.88083, 349.71042, 349.53925, 349.3675, 349.19525, 349.02237, 348.8487, 348.7615, 348.58633, 348.4099, 348.232, 348.0523, 347.87067, 347.68716, 347.50204, 347.31558, 347.12802, 346.92142, 346.7344, 346.5492, 346.3668, 346.1883, 346.0148, 345.84747, 345.68735, 345.53522, 345.39172, 345.25754, 345.13324, 345.019, 344.91495, 344.821, 344.73724, 344.6631, 344.59787, 344.54092, 344.49152, 344.46942, 344.43, 344.3962, 344.3674, 344.34283, 344.32196, 344.30417, 344.28894, 344.2756, 344.26346, 344.25177, 344.24585, 344.23355, 344.22025, 344.20566, 344.18954, 344.1716, 344.15182, 344.1303, 344.10715, 344.08237, 344.0562, 344.04266, 344.01474, 343.98593, 343.9565, 343.92685, 343.8974, 343.86853, 343.8405, 343.8134, 343.78717, 343.76184, 343.7373, 343.7132, 343.68918, 343.66486, 343.63974, 343.61304, 343.58398, 343.55176, 343.51575, 343.47543, 343.43045, 343.38037, 343.32486, 343.26385, 343.19727, 343.12506, 343.0473, 342.96426, 342.8763, 342.7838, 342.6871, 342.5868, 342.4834, 342.3775, 342.26956, 342.16, 342.04922, 341.9376, 341.8256, 341.71384, 341.603, 341.54816, 341.43988, 341.3337, 341.2298, 341.12817, 341.029, 340.93222, 340.83792, 340.74606, 340.65662, 340.61273, 340.5265, 340.44196, 340.3589, 340.27698, 340.1962, 340.11642, 340.03757, 339.9596, 339.8825, 339.80624, 339.76843, 339.69345, 339.61942, 339.5465, 339.4749, 339.40472, 339.33615, 339.26938, 339.20456, 339.17294, 339.11133, 339.0754, 339.01724, 338.96124, 338.90732, 338.85516, 338.80435, 338.7545, 338.70508, 338.65558, 338.60538, 338.55386, 338.50043, 338.44467, 338.38623, 338.3248, 338.26004, 338.19208, 338.12115, 338.04758, 337.97156, 337.8933, 337.813, 337.73077, 337.64688, 337.56183, 337.47614, 337.3905, 337.30548, 337.2219, 337.14047, 337.06207, 337.02423, 336.95163, 336.8833, 336.8195, 336.76038, 336.7059, 336.65552, 336.60852, 336.5643, 336.52222, 336.48163, 336.44193, 336.40244, 336.36282, 336.32297, 336.28293, 336.24268, 336.20255, 336.16336, 336.12595, 336.09125, 336.06015, 336.03354, 336.0124, 335.99765, 335.99005, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 335.94022, 335.8245, 335.7069, 335.5876, 335.4667, 335.34445, 335.22098, 335.09653, 334.9713, 334.84555, 334.7193, 334.59225, 334.46417, 334.3347, 334.2035, 334.07016, 333.9343, 333.79544, 333.65332, 333.5076, 333.3581, 333.20456, 333.04684, 332.88492, 332.7188, 332.54852, 332.37408, 332.19562, 332.0132, 331.827, 331.6372, 331.4442, 331.24854, 331.0506, 330.8508, 330.6493, 330.44623, 330.24173, 330.03598, 329.82928, 329.62195, 329.41428, 329.31042, 329.10284, 328.8958, 328.68967, 328.48474, 328.28125, 328.07925, 327.87888, 327.6802, 327.48328, 327.28802, 327.0945, 326.90268, 326.71255, 326.52423, 326.33774, 326.15317, 325.9707, 325.7906, 325.61313, 325.43854, 325.35233, 325.18204, 325.0145, 324.84952, 324.68692, 324.52628, 324.36713, 324.20905, 324.0517, 323.89508, 323.7392, 323.58417, 323.42996, 323.2766, 323.1242, 322.97272, 322.82224, 322.6728, 322.5245, 322.37738, 322.2315, 322.0867, 321.94275, 321.79953, 321.65692, 321.51486, 321.3734, 321.23264, 321.0925, 320.95316, 320.80096, 320.6637, 320.5276, 320.3927, 320.25916, 320.127, 319.9963, 319.86694, 319.7388, 319.6118, 319.48575, 319.36047, 319.23578, 319.11142, 318.98727, 318.86343, 318.73996, 318.617, 318.49466, 318.37314, 318.25266, 318.13342, 318.0743, 317.95706, 317.841, 317.72598, 317.61185, 317.49844, 317.38565, 317.27322, 317.16104, 317.04883, 316.93625, 316.82297, 316.7087, 316.59317, 316.4761, 316.35727, 316.23642, 316.1133, 315.98767, 315.85922, 315.72775, 315.59296, 315.4546, 315.31244, 315.16623, 315.016, 314.86185, 314.70395, 314.5425, 314.37762, 314.20947, 314.03818, 313.95142, 313.7758, 313.5977, 313.41745, 313.23547, 313.05212, 312.8678, 312.68286, 312.4977, 312.40518, 312.22037, 312.03616, 311.8529, 311.67087, 311.49026, 311.31122, 311.13388, 310.9583, 310.78464, 310.61276, 310.52753, 310.3584, 310.19098, 310.02484, 309.8595, 309.69455, 309.52945, 309.36377, 309.19702, 309.02872, 308.85843, 308.77246, 308.59866, 308.4222, 308.24283, 308.06033, 307.87457, 307.6854, 307.49268, 307.29626, 307.0758, 306.87122, 306.6626, 306.44995, 306.23343, 306.01324, 305.78952, 305.5626, 305.33286, 305.1007, 304.86655, 304.6307, 304.51227, 304.2745, 304.0359, 303.79666, 303.55713, 303.31754, 303.0781, 302.83896, 302.59998, 302.36093, 302.1216, 302.0018, 301.76187, 301.5215, 301.2807, 301.03943, 300.7977, 300.55554, 300.31293, 300.0699, 299.8264, 299.58237, 299.46017, 299.21527, 298.9699, 298.7245, 298.47946, 298.23532, 297.9924, 297.7507, 297.51016, 297.2707, 297.1513, 296.91293, 296.67456, 296.43564, 296.19553, 295.95374, 295.70978, 295.46323, 295.2136, 294.9607, 294.70456, 294.44516, 294.18253, 293.91678, 293.64816, 293.3769, 293.1033, 292.82773, 292.55078, 292.273, 291.995, 291.85614, 291.5792, 291.30402, 291.03152, 290.76245, 290.4973, 290.23663, 289.98083, 289.73035, 289.48505, 289.24493, 289.00986, 288.7797, 288.5541, 288.33267, 288.11502, 287.9008, 287.6898, 287.48178, 287.27658, 287.074, 286.87396, 286.6763, 286.481, 286.2879, 286.09705, 285.9084, 285.72195, 285.53772, 285.35553, 285.17526, 285.08582, 284.9082, 284.73215, 284.55756, 284.38422, 284.21204, 284.04095, 283.87097, 283.7021, 283.5344, 283.45105, 283.28558, 283.12213, 282.96106, 282.8028, 282.6476, 282.49573, 282.34744, 282.20297, 282.06235, 281.91217, 281.7798, 281.65125, 281.5262, 281.40433, 281.28522, 281.16846, 281.05365, 280.94046, 280.82846, 280.71722, 280.66177, 280.55078, 280.43933, 280.3269, 280.2132, 280.09784, 279.98056, 279.86115, 279.7397, 279.61655, 279.49216, 279.42963, 279.304, 279.17752, 279.05008, 278.9216, 278.7919, 278.66068, 278.52765, 278.39246, 278.25482, 278.11456, 278.04343, 277.89893, 277.7514, 277.6008, 277.44708, 277.29028, 277.1304, 276.96747, 276.80157, 276.6327, 276.46097, 276.37402, 276.19815, 276.01968, 275.8388, 275.6556, 275.4703, 275.28302, 275.0939, 274.9031, 274.71075, 274.51688, 274.4194, 274.22342, 274.02625, 273.82822, 273.62967, 273.43088, 273.2323, 273.03433, 272.83743, 272.642, 272.4485, 272.25717, 272.06845, 271.88263, 271.6999, 271.52032, 271.34406, 271.1711, 271.00134, 270.8344, 270.66995, 270.5076, 270.347, 270.1877, 270.02936, 269.87152, 269.71396, 269.5566, 269.39935, 269.2421, 269.0848, 269.00616, 268.84872, 268.6912, 268.5335, 268.37582, 268.2183, 268.06107, 267.90427, 267.748, 267.57666, 267.4215, 267.2669, 267.11282, 266.95923, 266.806, 266.65314, 266.50055, 266.34814, 266.1959, 266.04373, 265.96777, 265.81622, 265.6654, 265.51556, 265.36682, 265.2193, 265.07306, 264.9282, 264.78464, 264.6423, 264.501, 264.3607, 264.22137, 264.08322, 263.94644, 263.81122, 263.6775, 263.545, 263.41364, 263.2831, 263.15323, 263.08847, 262.95926, 262.83023, 262.7012, 262.57193, 262.44214, 262.31158, 262.18002, 262.0474, 261.91376, 261.84653, 261.71124, 261.5749, 261.43756, 261.29922, 261.16, 261.02008, 260.87973, 260.7393, 260.59906, 260.4594, 260.32077, 260.25198, 260.1157, 259.98138, 259.84897, 259.71832, 259.58926, 259.46164, 259.33533, 259.21027, 259.08627, 258.9633, 258.84128, 258.72018, 258.59998, 258.48056, 258.3617, 258.24307, 258.12436, 258.0053, 257.88574, 257.8257, 257.7051, 257.58356, 257.461, 257.33722, 257.2121, 257.08545, 256.95706, 256.8266, 256.6937, 256.5581, 256.41962, 256.34927, 256.20654, 256.06097, 255.91273, 255.76224, 255.60999, 255.45648, 255.30219, 255.1473, 254.99197, 254.8364, 254.68071, 254.52522, 254.37021, 254.21597, 254.06277, 253.9106, 253.75945, 253.60925, 253.46, 253.37088, 253.22295, 253.07571, 252.92911, 252.78325, 252.63849, 252.49512, 252.35345, 252.21367, 252.07579, 252.0076, 251.87268, 251.73972, 251.60844, 251.47859, 251.34984, 251.22192, 251.09464, 250.96782, 250.84126, 250.71481, 250.58826, 250.46143, 250.33415, 250.20624, 250.07756, 249.94798, 249.81737, 249.68564, 249.55289, 249.41924, 249.35213, 249.21738, 249.0821, 248.94655, 248.81093, 248.67545, 248.54044, 248.40631, 248.27348, 248.14236, 248.01303, 247.88528, 247.75894, 247.63379, 247.5096, 247.38615, 247.26318, 247.14049, 247.01793, 246.89554, 246.77333, 246.6513, 246.52962, 246.40848, 246.28815, 246.16884, 246.05067, 245.93369, 245.81789, 245.70326, 245.58977, 245.47722, 245.36548, 245.30986, 245.19904, 245.08864, 244.97852, 244.86853}
tdry =
  {28.2, 28.452778, 28.425447, 28.397804, 28.369694, 28.340958, 28.311445, 28.281, 28.249472, 28.216711, 28.182606, 28.147049, 28.109938, 28.071188, 28.030823, 27.988894, 27.945448, 27.900574, 27.854506, 27.807518, 27.75989, 27.711887, 27.663748, 27.615692, 27.56795, 27.520731, 27.474195, 27.428486, 27.383745, 27.340084, 27.297476, 27.255848, 27.215134, 27.175262, 27.136168, 27.097776, 27.060022, 27.022846, 26.986256, 26.950272, 26.91492, 26.880224, 26.846212, 26.812916, 26.780363, 26.748592, 26.717667, 26.687666, 26.658669, 26.630754, 26.604044, 26.578663, 26.554739, 26.532417, 26.511915, 26.49347, 26.477324, 26.463724, 26.452948, 26.445284, 26.440788, 26.440592, 26.444393, 26.452478, 26.46513, 26.48259, 26.504944, 26.53224, 26.564528, 26.601784, 26.643717, 26.689974, 26.740194, 26.79394, 26.850445, 26.908861, 26.968342, 27.028133, 27.087852, 27.147217, 27.20594, 27.263775, 27.320618, 27.376402, 27.431063, 27.484404, 27.535692, 27.584055, 27.62862, 27.668621, 27.703766, 27.733889, 27.758814, 27.778456, 27.793055, 27.802948, 27.808468, 27.80992, 27.807468, 27.801245, 27.791376, 27.778017, 27.76141, 27.741829, 27.71955, 27.694813, 27.667734, 27.638391, 27.606861, 27.57321, 27.537464, 27.499628, 27.459717, 27.417763, 27.37392, 27.328379, 27.28133, 27.232948, 27.18336, 27.13267, 27.080988, 27.028444, 26.975294, 26.921827, 26.86833, 26.8151, 26.762468, 26.710773, 26.660355, 26.611528, 26.564499, 26.519436, 26.476505, 26.43585, 26.397455, 26.361258, 26.327196, 26.295189, 26.26503, 26.23648, 26.2093, 26.183247, 26.158098, 26.13363, 26.109621, 26.085855, 26.062166, 26.0384, 26.014406, 25.990046, 25.965279, 25.940098, 25.914492, 25.88845, 25.861944, 25.834932, 25.80738, 25.779259, 25.75058, 25.718428, 25.688677, 25.658472, 25.627893, 25.597038, 25.566, 25.534864, 25.503695, 25.472544, 25.441467, 25.410505, 25.379631, 25.348803, 25.317978, 25.287117, 25.256191, 25.225178, 25.194052, 25.162786, 25.131342, 25.099676, 25.067743, 25.035484, 25.002779, 24.969484, 24.935455, 24.900553, 24.864634, 24.827562, 24.789196, 24.749414, 24.708164, 24.665417, 24.621147, 24.575354, 24.52817, 24.47977, 24.430334, 24.38007, 24.329374, 24.278696, 24.228485, 24.179163, 24.130991, 24.084188, 24.03897, 23.99555, 23.954107, 23.914808, 23.877825, 23.843285, 23.81109, 23.78108, 23.753094, 23.726952, 23.702417, 23.679234, 23.657145, 23.63591, 23.615385, 23.595453, 23.576002, 23.556944, 23.538322, 23.520231, 23.50276, 23.485989, 23.469923, 23.454548, 23.439844, 23.425774, 23.41219, 23.398901, 23.385721, 23.372467, 23.359016, 23.345259, 23.331085, 23.316397, 23.301146, 23.285297, 23.268826, 23.251705, 23.233965, 23.21565, 23.19681, 23.177477, 23.157654, 23.137316, 23.116446, 23.095032, 23.0731, 23.050697, 23.027868, 23.00466, 22.981146, 22.95741, 22.933537, 22.909601, 22.885656, 22.861746, 22.837908, 22.814182, 22.790604, 22.764875, 22.741705, 22.718775, 22.696108, 22.673721, 22.651634, 22.629862, 22.608381, 22.587168, 22.56619, 22.545422, 22.524818, 22.50434, 22.483942, 22.463596, 22.443354, 22.423292, 22.403486, 22.384014, 22.36496, 22.346409, 22.328453, 22.311161, 22.294537, 22.278559, 22.263206, 22.248417, 22.233917, 22.219358, 22.204401, 22.188738, 22.172295, 22.155066, 22.137045, 22.11826, 22.098879, 22.079128, 22.059233, 22.03942, 22.019926, 22.001005, 21.9829, 21.965853, 21.950037, 21.935614, 21.922747, 21.911602, 21.902412, 21.89543, 21.890903, 21.88905, 21.88988, 21.893328, 21.899332, 21.907803, 21.918495, 21.931112, 21.945358, 21.960934, 21.977562, 21.994967, 22.012875, 22.031004, 22.049057, 22.06672, 22.08368, 22.099651, 22.11448, 22.128063, 22.140303, 22.15111, 22.16046, 22.168362, 22.174822, 22.179857, 22.183558, 22.186047, 22.187445, 22.187868, 22.18742, 22.18619, 22.18427, 22.181736, 22.17851, 22.174461, 22.169456, 22.163353, 22.15593, 22.146935, 22.136114, 22.123247, 22.108303, 22.091333, 22.072388, 22.051521, 22.028786, 22.004236, 21.977926, 21.949883, 21.919903, 21.887691, 21.852953, 21.811491, 21.770649, 21.72666, 21.679388, 21.62875, 21.57497, 21.518373, 21.459288, 21.398045, 21.334995, 21.270506, 21.204939, 21.138638, 21.071829, 21.004694, 20.937424, 20.870222, 20.803417, 20.737381, 20.672483, 20.609056, 20.547218, 20.48701, 20.428469, 20.371603, 20.316225, 20.262075, 20.208899, 20.156437, 20.10444, 20.052668, 20.000872, 19.948835, 19.896488, 19.843813, 19.790794, 19.737452, 19.684006, 19.63076, 19.57801, 19.526072, 19.475336, 19.426228, 19.37917, 19.334549, 19.292522, 19.253155, 19.216515, 19.182653, 19.151522, 19.123035, 19.097103, 19.07361, 19.05224, 19.032597, 19.01428, 18.996895, 18.98003, 18.963272, 18.946205, 18.928436, 18.90973, 18.889917, 18.868822, 18.846275, 18.822123, 18.79622, 18.768423, 18.738585, 18.706553, 18.672173, 18.635294, 18.59576, 18.553425, 18.508137, 18.459747, 18.408112, 18.353138, 18.294752, 18.23288, 18.167461, 18.098526, 18.026146, 17.95039, 17.871347, 17.789255, 17.704416, 17.61713, 17.52773, 17.436785, 17.344965, 17.252945, 17.152271, 17.061787, 16.972736, 16.885548, 16.800598, 16.717945, 16.637526, 16.559282, 16.483149, 16.40899, 16.336658, 16.265997, 16.196861, 16.129137, 16.062729, 15.997536, 15.933457, 15.8703985, 15.808261, 15.746947, 15.686363, 15.626424, 15.567049, 15.508159, 15.449671, 15.391487, 15.333505, 15.27562, 15.217736, 15.1597805, 15.101693, 15.043416, 14.984893, 14.926106, 14.86705, 14.80772, 14.748108, 14.688179, 14.627892, 14.567202, 14.506067, 14.444456, 14.3823395, 14.319687, 14.256473, 14.1926985, 14.128372, 14.063504, 13.998109, 13.932221, 13.865889, 13.799157, 13.732078, 13.664722, 13.597176, 13.529523, 13.4618435, 13.394188, 13.326592, 13.259092, 13.191721, 13.124468, 13.057305, 12.990206, 12.923146, 12.856137, 12.789203, 12.722366, 12.655655, 12.589102, 12.522745, 12.456622, 12.390773, 12.32525, 12.260112, 12.19542, 12.131247, 12.067769, 12.005213, 11.943804, 11.8837805, 11.82547, 11.769239, 11.715459, 11.66449, 11.616632, 11.57216, 11.531341, 11.494434, 11.461585, 11.432883, 11.408419, 11.388262, 11.372326, 11.360443, 11.352446, 11.34813, 11.346985, 11.348339, 11.351523, 11.3558655, 11.360686, 11.365302, 11.369028, 11.371201, 11.371345, 11.369081, 11.364029, 11.355842, 11.344425, 11.329823, 11.312079, 11.289013, 11.265048, 11.238529, 11.209743, 11.178967, 11.14642, 11.1122875, 11.076758, 11.040002, 11.002046, 10.962861, 10.922417, 10.880692, 10.837718, 10.793554, 10.748256, 10.701891, 10.6546, 10.606553, 10.557923, 10.5088825, 10.459606, 10.410272, 10.361056, 10.312138, 10.2637, 10.215928, 10.169011, 10.123126, 10.078391, 10.034901, 9.992745, 9.95201, 9.912731, 9.874918, 9.838582, 9.803728, 9.770305, 9.738236, 9.707447, 9.677855, 9.649345, 9.621791, 9.595061, 9.569025, 9.543561, 9.518548, 9.493864, 9.46939, 9.445009, 9.42061, 9.396081, 9.371309, 9.346203, 9.320679, 9.294654, 9.268046, 9.2408085, 9.212907, 9.184307, 9.154978, 9.124886, 9.094001, 9.062291, 9.029724, 8.996244, 8.961785, 8.92628, 8.889666, 8.85191, 8.813, 8.772921, 8.731664, 8.689258, 8.645756, 8.601212, 8.555679, 8.509238, 8.461985, 8.414009, 8.365407, 8.316262, 8.266654, 8.216663, 8.166369, 8.115879, 8.065308, 8.0147705, 7.9643793, 7.9141827, 7.8641944, 7.814428, 7.75996, 7.710737, 7.661846, 7.6133375, 7.565257, 7.5176015, 7.4703474, 7.4234715, 7.376951, 7.3307705, 7.2849174, 7.239378, 7.194141, 7.149195, 7.104532, 7.0601416, 7.0160027, 6.9719977, 6.927966, 6.883746, 6.839171, 6.7940283, 6.748086, 6.701111, 6.6529107, 6.6036215, 6.5535355, 6.5029473, 6.4521484, 6.4014115, 6.3510003, 6.301179, 6.2521873, 6.204064, 6.1567492, 6.1101832, 6.0642824, 6.0187764, 5.9733, 5.9274874, 5.8809867, 5.833574, 5.785089, 5.7353725, 5.684271, 5.631682, 5.5775304, 5.5217404, 5.464266, 5.4053216, 5.3452587, 5.2844296, 5.2231884, 5.161908, 5.1009703, 5.040757, 4.98164, 4.9238877, 4.8677154, 4.813337, 4.7609625, 4.710766, 4.662901, 4.617521, 4.57477, 4.534701, 4.497316, 4.462616, 4.43056, 4.40069, 4.372314, 4.3447366, 4.3172836, 4.289495, 4.261033, 4.231562, 4.2007885, 4.1688576, 4.13617, 4.1031294, 4.070138, 4.0375957, 4.005898, 3.975441, 3.9465933, 3.91943, 3.8938518, 3.8697555, 3.847026, 3.8254068, 3.8045547, 3.7841265, 3.7637973, 3.7434485, 3.7230904, 3.702734, 3.6823921, 3.6620936, 3.6418774, 3.621783, 3.6018515, 3.5821555, 3.5608706, 3.5419662, 3.5235717, 3.5056984, 3.4883218, 3.471417, 3.454962, 3.438961, 3.42343, 3.408385, 3.3938422, 3.3798199, 3.3663366, 3.3534105, 3.341055, 3.3292298, 3.3178697, 3.306908, 3.296281, 3.2859492, 3.275884, 3.2660575, 3.2564461, 3.2470653, 3.2379506, 3.2291386, 3.2206638, 3.212549, 3.2048101, 3.1974633, 3.1905239, 3.1839967, 3.177882, 3.1721797, 3.1668875, 3.1619802, 3.1574194, 3.1531675, 3.1491842, 3.1454134, 3.141789, 3.138245, 3.1347146, 3.1311204, 3.127379, 3.1234071, 3.1191216, 3.1144378, 3.1092715, 3.1035373, 3.097158, 3.0901287, 3.0863822, 3.07845, 3.0699642, 3.060968, 3.0515158, 3.0416634, 3.0314658, 3.0209668, 3.010182, 2.9991233, 2.9878032, 2.976224, 2.9643662, 2.9522076, 2.9397259, 2.9268866, 2.9136264, 2.8998787, 2.8855765, 2.8706546, 2.8550544, 2.838718, 2.8215873, 2.8036072, 2.7847292, 2.7649066, 2.7440922, 2.7222683, 2.6994917, 2.67583, 2.65135, 2.626108, 2.6001282, 2.5734317, 2.5460389, 2.517974, 2.489271, 2.4599652, 2.4300926, 2.399695, 2.368832, 2.337566, 2.3059585, 2.2740734, 2.2419777, 2.2097385, 2.1774232, 2.1451063, 2.1128783, 2.080834, 2.0459092, 2.0145674, 1.9837455, 1.9535733, 1.9241818, 1.8957065, 1.8682956, 1.8420981, 1.8172635, 1.7939407, 1.7722784, 1.7524252, 1.7345295, 1.7186666, 1.7047566, 1.6927003, 1.6823972, 1.6736556, 1.6660854, 1.65927, 1.6527936, 1.6462479, 1.6392423, 1.6313889, 1.6222999, 1.6116568, 1.5992953, 1.5850717, 1.5688432, 1.5505437, 1.5302811, 1.5081873, 1.4843947, 1.4590583, 1.4323864, 1.4045948, 1.3758992, 1.3465259, 1.3167269, 1.2867576, 1.2568729, 1.2272884, 1.1981256, 1.1694921, 1.1414956, 1.1142083, 1.0876176, 1.0616983, 1.0364249, 1.0116976, 0.9872354, 0.96272963, 0.937872, 0.9123791, 0.8860299, 0.8586128, 0.8299163, 0.7998238, 0.7684569, 0.7359743, 0.70253485, 0.66831994, 0.63356906, 0.5985309, 0.563454, 0.5285552, 0.49396965, 0.45981887, 0.42622456, 0.39327943, 0.36099982, 0.32938966, 0.29845273, 0.2681634, 0.23841706, 0.2090958, 0.18008189, 0.15126093, 0.122528024, 0.093779825, 0.06491301, 0.035838906, 0.0065093343, -0.023116928, -0.05308109, -0.083418205, -0.114145935, -0.14527893, -0.17683187, -0.20882642, -0.24130443, -0.27431127, -0.30789232, -0.34207192, -0.3768134, -0.4120691, -0.4477913, -0.4839223, -0.5203746, -0.5570553, -0.5938716, -0.63076794, -0.67151517, -0.70878905, -0.7463631, -0.7843025, -0.82264346, -0.86141825, -0.900659, -0.9403781, -0.9805415, -1.0211086, -1.0620393, -1.1033162, -1.1449779, -1.1870707, -1.2296407, -1.2727071, -1.3162245, -1.3601379, -1.4043925, -1.448898, -1.4934789, -1.537947, -1.5821142, -1.6257603, -1.6685873, -1.7102855, -1.7505451, -1.7890847, -1.8256928, -1.8601692, -1.8923135, -1.921951, -1.9489716, -1.9732751, -1.9947615, -2.0133407, -2.0289488, -2.0415256, -2.0510116, -2.0573595, -2.060558, -2.0609746, -2.0594375, -2.0547462, -2.047038, -2.0365438, -2.023496, -2.0081296, -1.9907221, -1.9715788, -1.9510064, -1.9293118, -1.9068091, -1.8838178, -1.8606576, -1.8376544, -1.8152252, -1.793853, -1.7740222, -1.7562143, -1.7408695, -1.7283981, -1.7192096, -1.7136977, -1.7120366, -1.7142352, -1.7202986, -1.7302239, -1.7438889, -1.7610809, -1.7815852, -1.8051847, -1.8316284, -1.8606393, -1.8919395, -1.925252, -1.9603059, -1.9968367, -2.0345788, -2.0732667, -2.1126165, -2.152331, -2.1921122, -2.2316632, -2.27071, -2.3089948, -2.3462613, -2.3822567, -2.4168031, -2.4497817, -2.4810762, -2.510575, -2.5382488, -2.5641367, -2.58828, -2.6107244, -2.631589, -2.6510541, -2.669303, -2.6865168, -2.7028532, -2.7184503, -2.7334456, -2.7479787, -2.7622302, -2.7764156, -2.7907522, -2.8054583, -2.8207862, -2.8370168, -2.854432, -2.8733091, -2.8938317, -2.918428, -2.9427326, -2.9689846, -2.9971983, -3.0273337, -3.0593505, -3.093204, -3.1288066, -3.16604, -3.2047849, -3.2449214, -3.2863195, -3.328841, -3.3723483, -3.4167056, -3.461812, -3.5075912, -3.553967, -3.6008651, -3.648232, -3.6960287, -3.7200763, -3.7684462, -3.8171494, -3.8661442, -3.915388, -3.964839, -4.0144567, -4.064206, -4.114054, -4.1639667, -4.2139096, -4.263848, -4.313745, -4.363566, -4.4132657, -4.4627748, -4.5120196, -4.5609255, -4.6094255, -4.6574707, -4.705017, -4.75202, -4.7984476, -4.8443108, -4.8896265, -4.9344125, -4.9786963, -5.022538, -5.066004, -5.1091585, -5.152065, -5.1947694, -5.237317, -5.2797523, -5.3221, -5.3643217, -5.406365, -5.448178, -5.489708, -5.530897, -5.5716867, -5.612018, -5.6518517, -5.691211, -5.7301354, -5.768662, -5.806836, -5.844732, -5.882429, -5.9200063, -5.9575295, -5.995012, -6.0324574, -6.069868, -6.107243, -6.1445646, -6.1818123, -6.2189646, -6.256005, -6.292926, -6.3297253, -6.3663993, -6.4029408, -6.4393253, -6.475528, -6.51152, -6.5472713, -6.5827346, -6.6178594, -6.652595, -6.6868925, -6.7207108, -6.7540107, -6.786752, -6.8189197, -6.8505826, -6.881831, -6.9127564, -6.943468, -6.974148, -7.0049953, -7.03621, -7.055195, -7.0873513, -7.120242, -7.153972, -7.1886415, -7.2242894, -7.2609043, -7.298476, -7.336993, -7.376446, -7.416826, -7.4581246, -7.5003304, -7.5433674, -7.587109, -7.6314287, -7.6761947, -7.7212253, -7.766295, -7.811178, -7.8556523, -7.899537, -7.9426885, -7.9849634, -8.026223, -8.066408, -8.105519, -8.143564, -8.180546, -8.216465, -8.251316, -8.285094, -8.317796, -8.3494215, -8.379983, -8.409489, -8.43795, -8.465411, -8.491946, -8.517628, -8.542527, -8.566678, -8.590077, -8.612721, -8.634606, -8.655687, -8.675888, -8.695129, -8.713336, -8.730495, -8.746652, -8.761849, -8.776138, -8.7896385, -8.802531, -8.815002, -8.82724, -8.839499, -8.852098, -8.865355, -8.879584, -8.895012, -8.9117775, -8.930018, -8.949864, -8.971305, -8.994192, -9.018374, -9.043699, -9.0700035, -9.097114, -9.124858, -9.153064, -9.181572, -9.210238, -9.238919, -9.267469, -9.295727, -9.323511, -9.350644, -9.376945, -9.402269, -9.41453, -9.43818, -9.460575, -9.481635, -9.501394, -9.519917, -9.537268, -9.553536, -9.568929, -9.5836735, -9.599424, -9.613577, -9.627852, -9.642531, -9.657891, -9.674189, -9.691603, -9.7103, -9.730446, -9.752178, -9.775558, -9.800628, -9.827428, -9.855981, -9.886236, -9.918127, -9.9515915, -9.986558, -10.022944, -10.060667, -10.099638, -10.139781, -10.18104, -10.223365, -10.2667055, -10.311026, -10.356334, -10.40265, -10.449991, -10.498404, -10.548023, -10.599005, -10.6515045, -10.705633, -10.761346, -10.81856, -10.877195, -10.937117, -10.997993, -11.059452, -11.121119, -11.182619, -11.243587, -11.3036585, -11.362468, -11.419678, -11.475053, -11.528382, -11.579454, -11.628113, -11.674403, -11.696691, -11.73961, -11.780405, -11.81927, -11.85649, -11.892353, -11.927146, -11.961097, -11.994378, -12.027158, -12.059603, -12.091778, -12.12365, -12.155179, -12.186327, -12.216994, -12.247027, -12.276269, -12.30456, -12.331725, -12.357569, -12.381897, -12.404516, -12.425302, -12.444196, -12.461145, -12.476103, -12.489137, -12.500439, -12.510208, -12.518645, -12.525982, -12.532486, -12.538429, -12.54408, -12.54971, -12.555593, -12.561998, -12.5692005, -12.577444, -12.586949, -12.597931, -12.604044, -12.617617, -12.633002, -12.6502, -12.66921, -12.690018, -12.712535, -12.736655, -12.762269, -12.789274, -12.820477, -12.850109, -12.880859, -12.912653, -12.945465, -12.979277, -13.014072, -13.049842, -13.086602, -13.124373, -13.1631775, -13.203047, -13.244046, -13.286252, -13.32974, -13.374572, -13.420763, -13.468318, -13.51724, -13.567527, -13.619154, -13.6720915, -13.726311, -13.781777, -13.838448, -13.896276, -13.955215, -14.015211, -14.07618, -14.138031, -14.200671, -14.264007, -14.327926, -14.392313, -14.457054, -14.522024, -14.587061, -14.651991, -14.716641, -14.780828, -14.844317, -14.906859, -14.968209, -15.028144, -15.086556, -15.143367, -15.198495, -15.251886, -15.303585, -15.353664, -15.402196, -15.449265, -15.49501, -15.539588, -15.583152, -15.625859, -15.667873, -15.709363, -15.750493, -15.791412, -15.832191, -15.872875, -15.913511, -15.954142, -15.994782, -16.035442, -16.076132, -16.116867, -16.157701, -16.198698, -16.239918, -16.281404, -16.323107, -16.364944, -16.406837, -16.448706, -16.490448, -16.531961, -16.57314, -16.613886, -16.65414, -16.693855, -16.732975, -16.771461, -16.809292, -16.846458, -16.88295, -16.918758, -16.953876, -16.988304, -17.022038, -17.055077, -17.071344, -17.103401, -17.134846, -17.16572, -17.196081, -17.22602, -17.255629, -17.284998, -17.314201, -17.343294, -17.375233, -17.404266, -17.433353, -17.46255, -17.491907, -17.52148, -17.551304, -17.581402, -17.611792, -17.642494, -17.673508, -17.70481, -17.736372, -17.768173, -17.800224, -17.832573, -17.865263, -17.898346, -17.931826, -17.965664, -17.999823, -18.034266, -18.068956, -18.103867, -18.138966, -18.174227, -18.209639, -18.245213, -18.28096, -18.316895, -18.353016, -18.389318, -18.42579, -18.462427, -18.499231, -18.53623, -18.573446, -18.610905, -18.648628, -18.686634, -18.724947, -18.763584, -18.802538, -18.84177, -18.881243, -18.920916, -18.960747, -19.000704, -19.040749, -19.080841, -19.120918, -19.160875, -19.20061, -19.240015, -19.278936, -19.317156, -19.354454, -19.3906, -19.42509, -19.45709, -19.48574, -19.51021, -19.53036, -19.546911, -19.560637, -19.572304, -19.582682, -19.592525, -19.602598, -19.613651, -19.626211, -19.640518, -19.6484, -19.66575, -19.685383, -19.70731, -19.731497, -19.757904, -19.786482, -19.817104, -19.849623, -19.88389, -19.919754, -19.957048, -19.995598, -20.03523, -20.07578, -20.117138, -20.159204, -20.201885, -20.24509, -20.288757, -20.332842, -20.377295, -20.422064, -20.467093, -20.512321, -20.557692, -20.60314, -20.648619, -20.69408, -20.739477, -20.784752, -20.829803, -20.874512, -20.918755, -20.96242, -21.005426, -21.047714, -21.08922, -21.129889, -21.169748, -21.20885, -21.251059, -21.288746, -21.325808, -21.362251, -21.398088, -21.433338, -21.468033, -21.50222, -21.535942, -21.56925, -21.602224, -21.634956, -21.667536, -21.70005, -21.732574, -21.765177, -21.797922, -21.830872, -21.864038, -21.897419, -21.931015, -21.964823, -21.99883, -22.03303, -22.067404, -22.101944, -22.13666, -22.17156, -22.20666, -22.241966, -22.277458, -22.313112, -22.3489, -22.384796, -22.420752, -22.456724, -22.492662, -22.528524, -22.564312, -22.600039, -22.635714, -22.67135, -22.706963, -22.74256, -22.778154, -22.813759, -22.849392, -22.885075, -22.920828, -22.956675, -22.992634, -23.02873, -23.064991, -23.10143, -23.138046, -23.17483, -23.211765, -23.248846, -23.28608, -23.32348, -23.361069, -23.39885, -23.436808, -23.474913, -23.513136, -23.55144, -23.589733, -23.627907, -23.665848, -23.703447, -23.740608, -23.777239, -23.813248, -23.848547, -23.883095, -23.916866, -23.949835, -23.981983, -24.013311, -24.043837, -24.073574, -24.102545, -24.13084, -24.15857, -24.185844, -24.212788, -24.239594, -24.266485, -24.293684, -24.32141, -24.349854, -24.379192, -24.409609, -24.441284, -24.474419, -24.509224, -24.545912, -24.584673, -24.625599, -24.668736, -24.714125, -24.761797, -24.816736, -24.868776, -24.922642, -24.978151, -25.035069, -25.093132, -25.152082, -25.211655, -25.271576, -25.331568, -25.391348, -25.450636, -25.509132, -25.566534, -25.62254, -25.676859, -25.729273, -25.779598, -25.82764, -25.873232, -25.916304, -25.956827, -25.99477, -26.030128, -26.06304, -26.093693, -26.12228, -26.149002, -26.17414, -26.198008, -26.220911, -26.243147, -26.264936, -26.286469, -26.307936, -26.329521, -26.351381, -26.373652, -26.396479, -26.419987, -26.444227, -26.469221, -26.494987, -26.521542, -26.548838, -26.57681, -26.605396, -26.634535, -26.664213, -26.69444, -26.72522, -26.756548, -26.788355, -26.820553, -26.853045, -26.885738, -26.918518, -26.951262, -26.983847, -27.01616, -27.048128, -27.079704, -27.110832, -27.141474, -27.171635, -27.20135, -27.23065, -27.259571, -27.288185, -27.316568, -27.344803, -27.372969, -27.401152, -27.415274, -27.443634, -27.472216, -27.501076, -27.530216, -27.559643, -27.589354, -27.619368, -27.649717, -27.68044, -27.695953, -27.727297, -27.759026, -27.791082, -27.82341, -27.855944, -27.888597, -27.921274, -27.953876, -27.986305, -28.02162, -28.05325, -28.084278, -28.114563, -28.143927, -28.172178, -28.19913, -28.224594, -28.248415, -28.270435, -28.290504, -28.308477, -28.324278, -28.33785, -28.34914, -28.358112, -28.364862, -28.369532, -28.372263, -28.373215, -28.3731, -28.37188, -28.369581, -28.366503, -28.362976, -28.359383, -28.35611, -28.353546, -28.352098, -28.352205, -28.354313, -28.356253, -28.362152, -28.370882, -28.382568, -28.397333, -28.415272, -28.436266, -28.460125, -28.486654, -28.515636, -28.54669, -28.562857, -28.596191, -28.63049, -28.665276, -28.700024, -28.734198, -28.767271, -28.798744, -28.828178, -28.855137, -28.879187, -28.899933, -28.917048, -28.930214, -28.939104, -28.943247, -28.941925, -28.9344, -28.919943, -28.898533, -28.871298, -28.839474, -28.8043, -28.767132, -28.729511, -28.693005, -28.65917, -28.629135, -28.603302, -28.582003, -28.565565, -28.55414, -28.547564, -28.54564, -28.54818, -28.554909, -28.565416, -28.579287, -28.596092, -28.615395, -28.636702, -28.659523, -28.671349, -28.695534, -28.720133, -28.74482, -28.769264, -28.793154, -28.81629, -28.838524, -28.859713, -28.879717, -28.889248, -28.907335, -28.924082, -28.93944, -28.953386, -28.96595, -28.977169, -28.987076, -28.995708, -29.0031, -29.009283, -29.011932, -29.016365, -29.01968, -29.021915, -29.023108, -29.023298, -29.022514, -29.02078, -29.018122, -29.016453, -29.012447, -29.009619, -29.004208, -28.997934, -28.990826, -28.983019, -28.974695, -28.966038, -28.957237, -28.948566, -28.940327, -28.93282, -28.926325, -28.92094, -28.916689, -28.913597, -28.911678, -28.91086, -28.911037, -28.912104, -28.913944, -28.916424, -28.919386, -28.922678, -28.92614, -28.929558, -28.932692, -28.935305, -28.937157, -28.937996, -28.937563, -28.935604, -28.933973, -28.929314, -28.922749, -28.91422, -28.90368, -28.891153, -28.876808, -28.860825, -28.84339, -28.82474, -28.805212, -28.785152, -28.76491, -28.744852, -28.725393, -28.706951, -28.689936, -28.674683, -28.661367, -28.65015, -28.641193, -28.634523, -28.629929, -28.627167, -28.626001, -28.626076, -28.626831, -28.627686, -28.628056, -28.62746, -28.625612, -28.62224, -28.617073, -28.609966, -28.601004, -28.590296, -28.57795, -28.564133, -28.549107, -28.533154, -28.516548, -28.508085, -28.490973, -28.473795, -28.456766, -28.440094, -28.423922, -28.40835, -28.393486, -28.379421, -28.366133, -28.353527, -28.34152, -28.330015, -28.31886, -28.307869, -28.296865, -28.285662, -28.274061, -28.261864, -28.248865, -28.233423, -28.21831, -28.202213, -28.18518, -28.167263, -28.148575, -28.129265, -28.109474, -28.089346, -28.069, -28.04855, -28.028103, -28.007767, -27.9876, -27.967646, -27.947945, -27.928532, -27.909409, -27.890566, -27.871986, -27.853666, -27.835653, -27.826784, -27.809364, -27.792433, -27.77604, -27.760204, -27.744946, -27.730278, -27.71621, -27.70273, -27.689833, -27.677505, -27.665724, -27.654448, -27.643631, -27.633228, -27.623152, -27.613237, -27.603317, -27.59322, -27.582838, -27.57218, -27.561272, -27.550133, -27.538826, -27.527494, -27.516283, -27.505342, -27.494797, -27.484737, -27.475248, -27.466412, -27.458292, -27.450907, -27.444271, -27.4384, -27.433323, -27.429104, -27.425812, -27.423512, -27.422277, -27.422192, -27.423336, -27.424398, -27.427544, -27.432085, -27.43805, -27.445461, -27.45433, -27.464573, -27.476038, -27.48858, -27.502018, -27.51582, -27.52926, -27.541615, -27.552177, -27.5605, -27.566265, -27.569162, -27.56895, -27.5661, -27.561491, -27.556005, -27.550491, -27.545414, -27.541012, -27.537527, -27.535185, -27.534071, -27.534187, -27.53554, -27.53812, -27.54187, -27.546688, -27.552475, -27.559128, -27.56649, -27.574375, -27.582602, -27.590982, -27.599325, -27.608229, -27.615866, -27.622871, -27.629097, -27.634413, -27.638687, -27.6418, -27.643682, -27.644302, -27.64362, -27.641603, -27.638287, -27.636156, -27.630985, -27.624653, -27.617357, -27.609573, -27.601803, -27.594551, -27.588457, -27.584421, -27.583368, -27.586227, -27.593792, -27.6066, -27.625158, -27.649973, -27.681013, -27.717201, -27.757332, -27.800209, -27.844837, -27.890636, -27.937075, -27.983622, -28.029854, -28.075556, -28.12054, -28.164618, -28.207668, -28.24971, -28.29078, -28.33091, -28.370155, -28.408598, -28.44633, -28.483438, -28.520023, -28.556202, -28.592096, -28.627827, -28.66351, -28.699257, -28.735182, -28.771393, -28.808004, -28.845135, -28.882904, -28.921432, -28.960825, -29.001162, -29.042513, -29.084951, -29.106592, -29.15065, -29.19564, -29.241438, -29.28791, -29.334923, -29.382332, -29.42999, -29.477762, -29.525547, -29.573277, -29.62088, -29.66829, -29.71545, -29.76232, -29.808851, -29.855005, -29.900757, -29.946095, -29.991007, -30.03548, -30.057543, -30.101282, -30.144468, -30.187046, -30.228964, -30.270166, -30.310606, -30.350227, -30.388975, -30.426771, -30.463543, -30.499212, -30.53373, -30.567118, -30.599403, -30.630617, -30.660809, -30.690077, -30.718525, -30.746264, -30.773384, -30.799969, -30.82609, -30.851818, -30.877207, -30.90224, -30.9269, -30.951164, -30.975002, -30.998371, -31.023483, -31.045725, -31.067383, -31.088495, -31.109098, -31.129236, -31.148964, -31.168365, -31.18753, -31.20655, -31.225494, -31.244398, -31.263287, -31.28219, -31.301126, -31.320086, -31.33906, -31.358038, -31.376997, -31.395887, -31.41466, -31.43326, -31.442486, -31.460802, -31.478975, -31.497047, -31.515059, -31.533072, -31.551157, -31.569386, -31.587828, -31.606565, -31.62568, -31.645264, -31.66539, -31.68611, -31.707445, -31.729418, -31.752056, -31.775377, -31.799408, -31.824167, -31.849682, -31.875969, -31.903055, -31.930964, -31.959705, -31.989197, -32.019287, -32.04982, -32.080654, -32.111683, -32.142838, -32.17404, -32.18964, -32.2208, -32.251904, -32.282936, -32.313892, -32.344776, -32.375656, -32.406605, -32.437687, -32.45331, -32.48479, -32.516735, -32.549297, -32.58263, -32.616817, -32.6519, -32.68792, -32.7249, -32.762844, -32.801704, -32.82147, -32.86164, -32.90267, -32.944656, -32.98771, -33.031937, -33.077385, -33.12391, -33.171326, -33.219467, -33.268105, -33.292503, -33.341236, -33.389572, -33.43714, -33.483475, -33.528027, -33.570255, -33.609634, -33.64592, -33.682224, -33.711914, -33.7385, -33.7627, -33.785656, -33.808506, -33.832336, -33.85769, -33.884777, -33.913815, -33.94499, -33.978333, -33.995796, -34.032257, -34.070705, -34.111015, -34.152927, -34.196167, -34.24046, -34.285587, -34.331467, -34.37803, -34.42521, -34.449017, -34.49709, -34.545807, -34.595222, -34.645374, -34.6963, -34.748016, -34.800537, -34.85388, -34.90806, -34.96305, -34.990852, -35.04706, -35.104042, -35.161694, -35.21991, -35.27857, -35.337593, -35.396976, -35.456726, -35.516846, -35.547054, -35.607887, -35.669445, -35.731937, -35.79557, -35.860405, -35.926407, -35.99354, -36.061768, -36.130898, -36.20067, -36.2708, -36.341, -36.410675, -36.47905, -36.545326, -36.608738, -36.66891, -36.72574, -36.779125, -36.828995, -36.8527, -36.898033, -36.941128, -36.982605, -37.022972, -37.062347, -37.10078, -37.13833, -37.175045, -37.210968, -37.246143, -37.280613, -37.314407, -37.34752, -37.379932, -37.411636, -37.442623, -37.472916, -37.502544, -37.53154, -37.559944, -37.58786, -37.6154, -37.642666, -37.66978, -37.696857, -37.724022, -37.751392, -37.779114, -37.807365, -37.836346, -37.85117, -37.881603, -37.91316, -37.945866, -37.97976, -38.01486, -38.05111, -38.088394, -38.12659, -38.16557, -38.1853, -38.225094, -38.265144, -38.305218, -38.3451, -38.384617, -38.42361, -38.461914, -38.499382, -38.5359, -38.57485, -38.60903, -38.64196, -38.673588, -38.703888, -38.732826, -38.76038, -38.786575, -38.811443, -38.835014, -38.85734, -38.868073, -38.888744, -38.908466, -38.927357, -38.945538, -38.963135, -38.980263, -38.997044, -39.013508, -39.02963, -39.045376, -39.0531, -39.068233, -39.082912, -39.097103, -39.110764, -39.12386, -39.136333, -39.14814, -39.159218, -39.169533, -39.179096, -39.1836, -39.19207, -39.19984, -39.207027, -39.21382, -39.220417, -39.227, -39.233845, -39.241253, -39.249542, -39.259026, -39.264282, -39.27591, -39.28914, -39.304096, -39.32087, -39.33942, -39.35968, -39.38158, -39.405064, -39.430088, -39.456615, -39.470432, -39.499153, -39.529297, -39.560852, -39.593803, -39.62813, -39.66383, -39.700874, -39.739254, -39.778954, -39.81992, -39.86208, -39.905354, -39.949665, -39.99489, -40.040874, -40.087463, -40.1345, -40.181843, -40.22937, -40.276943, -40.324444, -40.37169, -40.418476, -40.46459, -40.509808, -40.553894, -40.596573, -40.637558, -40.67659, -40.71354, -40.73123, -40.765064, -40.79683, -40.826565, -40.85444, -40.88064, -40.90536, -40.928802, -40.951202, -40.974926, -40.995926, -41.01662, -41.037205, -41.057873, -41.07881, -41.100174, -41.122013, -41.144356, -41.16724, -41.190674, -41.20258, -41.226715, -41.25123, -41.276047, -41.301117, -41.326412, -41.35189, -41.37753, -41.403336, -41.429363, -41.455654, -41.482258, -41.509197, -41.53648, -41.564117, -41.592113, -41.620464, -41.649147, -41.678146, -41.707436, -41.736977, -41.751823, -41.78162, -41.811504, -41.841423, -41.871326, -41.90118, -41.93094, -41.96056, -41.99001, -42.019257, -42.03379, -42.062656, -42.091236, -42.119503, -42.147434, -42.17501, -42.202156, -42.228775, -42.25476, -42.28001, -42.30447, -42.328117, -42.339626, -42.362007, -42.38355, -42.404377, -42.424637, -42.444473, -42.464016, -42.483356, -42.502575, -42.521744, -42.540936, -42.560192, -42.579544, -42.59903, -42.618668, -42.638485, -42.65849, -42.678696, -42.699104, -42.719685, -42.73003, -42.750797, -42.771637, -42.79256, -42.813614, -42.83484, -42.856293, -42.878105, -42.900494, -42.92367, -42.947853, -42.973125, -42.986164, -43.013016, -43.04088, -43.0697, -43.099327, -43.129593, -43.160328, -43.191395, -43.222755, -43.254406, -43.28634, -43.31854, -43.350986, -43.383644, -43.416485, -43.449482, -43.48264, -43.515953, -43.54944, -43.583096, -43.603367, -43.63727, -43.671314, -43.70548, -43.739754, -43.77412, -43.808563, -43.843075, -43.8777, -43.912537, -43.93007, -43.965412, -44.001213, -44.03758, -44.074604, -44.11239, -44.151005, -44.190434, -44.23064, -44.271584, -44.313236, -44.35556, -44.398533, -44.442127, -44.4863, -44.530975, -44.57606, -44.621468, -44.667107, -44.71287, -44.758648, -44.78151, -44.827106, -44.872417, -44.917286, -44.96155, -45.00505, -45.04762, -45.08906, -45.129196, -45.167835, -45.20482, -45.24002, -45.273296, -45.304516, -45.333366, -45.359386, -45.382114, -45.401108, -999.0, -45.428608, -45.438206, -45.445763, -45.451748, -45.456547, -45.460537, -45.464104, -45.46747, -45.470737, -45.473995, -45.477337, -45.48079, -45.484325, -45.487926, -45.48974, -45.493385, -45.497044, -45.500713, -45.504387}
dp =
  {16.152426, 15.808324, 15.752282, 15.696484, 15.641074, 15.586162, 15.531681, 15.477524, 15.42358, 15.369775, 15.316155, 15.262808, 15.209815, 15.157297, 15.105533, 15.054838, 15.005532, 14.957948, 14.912498, 14.869618, 14.829739, 14.793276, 14.760606, 14.732086, 14.708074, 14.688908, 14.67487, 14.6662245, 14.663229, 14.666071, 14.674637, 14.688724, 14.70813, 14.7325945, 14.761597, 14.794549, 14.830868, 14.869939, 14.910965, 14.95311, 14.995553, 15.037473, 15.07799, 15.116218, 15.151287, 15.182453, 15.209532, 15.232505, 15.251349, 15.266024, 15.276416, 15.282389, 15.283802, 15.280485, 15.272148, 15.258452, -999.0, 15.213694, 15.182553, 15.145953, 15.09975, 15.052567, 15.000284, 14.942625, 14.879288, 14.809971, 14.734443, 14.652472, 14.563795, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 12.992283, -999.0, -999.0, -999.0, 12.286886, 12.105842, 11.924498, 11.743115, 11.562018, 11.381545, 11.201911, 11.023297, 10.845893, 10.6699915, 10.496348, 10.325845, 10.159371, 9.99766, 9.840703, 9.688269, 9.540093, 9.395882, 9.255275, 9.117878, -999.0, 8.851085, 8.721347, 8.594184, 8.46972, 8.348067, 8.229294, 8.113451, 8.000586, 7.890769, -999.0, -999.0, 7.581795, 7.4864016, 7.3951197, 7.308094, 7.225463, 7.1473346, 7.0736804, 7.0044265, 6.9394937, 6.8787656, 6.821968, 6.7687764, 6.7188635, 6.6719265, 6.627789, 6.586314, 6.547364, 6.5108595, 6.4770107, 6.44612, 6.418489, 6.39438, 6.3738604, 6.3569307, 6.343592, 6.333789, 6.3271747, 6.3233104, 6.3217564, 6.3220406, 6.3235197, 6.3254967, 6.3272753, 6.328178, 6.3275943, 6.324941, 6.319638, 6.3112364, 6.3000093, 6.286474, 6.271145, 6.254523, 6.2370396, 6.217299, 6.1993318, 6.181766, 6.165022, 6.1495214, 6.1356845, 6.1238937, 6.1143737, 6.107305, 6.1028676, 6.101126, 6.1016626, 6.1039286, 6.1073804, 6.1114593, 6.115531, 6.1189446, 6.1210546, 6.121285, 6.1193514, 6.1150513, 6.108183, 6.0985727, 6.0861764, 6.0709867, 6.052993, 6.032156, 6.0083017, 5.9812183, 5.9506917, 5.9166436, 5.8796306, 5.8403935, 5.7996745, 5.7582235, 5.716833, 5.676309, 5.637454, 5.600971, 5.567087, 5.535882, 5.5074377, 5.4816647, 5.4576297, 5.434146, 5.4100337, 5.384226, 5.3561864, 5.3255444, 5.2919254, 5.2550654, 5.21527, 5.173026, 5.128818, 5.083093, 5.0361195, 4.9881053, 4.9392614, 4.889771, 4.8396564, 4.78889, 4.7374425, 4.6853065, 4.632584, 4.579413, 4.525933, 4.472282, 4.4185944, 4.3650045, 4.3116484, 4.2586665, 4.2062225, 4.154489, 4.103644, 4.053778, 4.0044823, 3.955169, 3.9052453, 3.8541267, 3.8012996, 3.7462716, 3.6885457, 3.6277516, 3.564287, 3.4988334, 3.4320805, 3.364769, 3.2979095, 3.232621, 3.1700354, 3.1112058, 3.0566542, 3.0067015, 2.9616654, 2.9218004, 2.8869932, 2.8569865, 2.831517, 2.810346, 2.7934117, 2.780719, 2.772269, 2.7681572, 2.7690878, 2.7770514, 2.7916012, 2.814042, 2.8452265, 2.8859732, 2.9370725, 2.9991949, 3.0725625, 3.1572437, 3.2532792, 3.3605978, 3.4786975, 3.606944, 3.7447004, 3.8912594, 4.0455694, 4.2065015, 4.3729677, -999.0, -999.0, 4.8951173, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 6.5843587, -999.0, -999.0, 6.9776177, -999.0, -999.0, -999.0, -999.0, -999.0, 7.556262, 7.6289935, -999.0, -999.0, -999.0, -999.0, -999.0, 7.9384103, -999.0, -999.0, -999.0, -999.0, 8.028375, 8.0282135, 8.021697, 8.008647, 7.988949, 7.962507, 7.929211, 7.889004, 7.842197, 7.7892385, 7.730581, 7.666748, 7.598661, 7.5274096, 7.454113, 7.379864, 7.3054147, 7.2313933, 7.158445, 7.0871587, 7.017702, 6.9500737, -999.0, -999.0, 6.7572594, 6.6946225, 6.631447, 6.5668964, 6.5002556, 6.430852, 6.357999, 6.2810726, 6.1999507, 6.1147203, 6.025471, 5.932347, 5.835841, 5.7366085, 5.635322, 5.5326695, 5.429309, 5.3258924, 5.2230835, 5.1215253, -999.0, -999.0, -999.0, 4.735538, 4.64612, 4.5607524, 4.4801507, 4.3978043, 4.329152, 4.2667456, 4.2108917, 4.1617866, 4.1190968, 4.082302, 4.050872, 4.0242586, 4.0018606, 3.9830618, 3.96725, -999.0, -999.0, 3.9305894, 3.9191263, 3.9066656, 3.8926399, -999.0, -999.0, -999.0, -999.0, 3.7837083, 3.752137, 3.716933, 3.6783483, 3.636761, 3.592544, 3.546086, 3.4978893, 3.4484963, 3.3984492, 3.3482533, 3.2981923, 3.2484682, 3.199283, 3.1508737, 3.1037006, 3.0583081, 3.0152388, 2.9750504, 2.9383974, 2.9059696, 2.878455, 2.8565018, 2.8405282, 2.83086, 2.8278165, 2.831689, 2.8425987, 2.8605988, 2.8857355, 2.9180038, 2.95709, 3.002554, 3.0539525, 3.110789, 3.1722412, 3.237359, 3.3052, 3.3748693, 3.4457433, 3.517313, 3.5890777, 3.6605332, 3.7311192, 3.800258, 3.867381, 3.931944, 3.993503, 4.0516605, 4.1060247, 4.156247, 4.2022576, 4.2441025, 4.2818246, 4.3154836, 4.3452964, 4.3715425, 4.3944955, 4.41446, 4.4320197, 4.447874, 4.4627085, 4.477137, 4.491341, 4.5053134, 4.519051, 4.5325656, 4.54594, 4.559299, 4.572782, -999.0, -999.0, 4.6172824, 4.6332607, 4.6503778, 4.6685834, 4.6877427, 4.707721, 4.7283115, 4.74886, 4.7685633, 4.786632, 4.802396, 4.8158193, 4.8270936, 4.836403, 4.8439445, 4.8500295, 4.8550053, 4.8592114, 4.8629823, 4.8666534, 4.870558, 4.8750215, 4.8803315, 4.886568, 4.8937316, 4.901819, 4.910807, 4.920544, 4.930834, 4.9414787, 4.9522386, 4.9625664, -999.0, -999.0, 4.984446, 4.986767, 4.9858594, 4.9813223, 4.9728117, 4.960339, 4.944058, 4.9241195, 4.900693, 4.874103, 4.844735, 4.8129716, 4.7792068, 4.7439604, 4.7078, 4.671289, 4.6349697, 4.5992565, 4.564509, 4.531082, 4.4992933, 4.4691935, 4.4407187, 4.413805, 4.3883843, 4.3643465, 4.341564, 4.3199096, 4.2992425, 4.27931, 4.2598124, 4.240453, 4.220957, 4.201185, 4.1810603, 4.1605062, 4.139462, 4.117969, 4.0961156, 4.07399, 4.0516424, 4.028825, 4.005153, 3.9802496, 3.9537215, 3.925026, 3.8935502, 3.8586843, 3.819828, 3.776461, 3.7280946, 3.674227, -999.0, -999.0, 3.4762235, 3.397853, -999.0, -999.0, -999.0, -999.0, -999.0, 2.8010728, 2.6814659, -999.0, -999.0, 2.288337, 2.1471145, 2.0019505, -999.0, -999.0, 1.5528661, -999.0, 1.2564162, 1.113554, 0.9760356, 0.8451881, 0.71050483, 0.59746414, 0.49410582, 0.40111262, 0.31903422, 0.24766214, 0.18644872, 0.13481161, 0.092111714, 0.057489205, 0.029983658, 0.0086226445, -0.0075453585, -0.01927983, -0.027257435, -0.032152902, -0.034624953, -0.035239626, -0.034518253, -0.032974172, -0.031081224, -0.029080808, -0.027110143, -0.02530166, -0.023709424, -0.021838699, -0.01895516, -0.014330734, -0.0072463555, 0.0029979388, 0.017087718, 0.03569816, 0.059435673, 0.08845746, 0.12271407, 0.16215298, 0.20663375, 0.2553495, 0.30719632, 0.36108992, 0.41597354, 0.4708573, 0.5247915, 0.5768437, 0.6261455, 0.6722295, -999.0, -999.0, -999.0, 0.818968, 0.8450922, 0.8666188, 0.8834306, 0.8959452, 0.9048396, 0.9107833, 0.91442114, 0.9162458, 0.91667235, 0.9161114, 0.9149239, 0.9130653, 0.9102852, 0.9063331, -999.0, -999.0, 0.88563436, 0.87554824, 0.86380213, 0.8505578, 0.8360778, 0.82062376, 0.80443025, 0.78750217, 0.76972234, 0.7509737, 0.73112184, 0.7098614, 0.68679607, -999.0, 0.6337245, 0.60347193, 0.57111466, 0.53699374, 0.5014575, 0.4649365, 0.42790666, 0.390843, 0.35421187, 0.31840822, 0.28378567, 0.2506957, 0.21645874, 0.18746671, 0.16057038, 0.13583072, 0.113261096, 0.092531286, 0.07316066, 0.05467126, 0.03662095, 0.01881117, 0.001153119, -0.016440887, -0.034039058, -0.05156622, -0.06888245, -0.08584865, -0.10233998, -0.11833379, -0.13385564, -0.14893256, -0.16358924, -0.1778235, -0.1916221, -0.20497431, -0.21785559, -0.23010948, -0.24151556, -0.25185266, -0.26093122, -0.2688201, -0.27571014, -0.2817875, -0.28723904, -0.2922983, -0.29722136, -0.30226237, -0.3076835, -0.31383124, -0.32109505, -0.3298648, -0.34050152, -0.3531176, -0.3677002, -0.38423726, -0.40272897, -0.4232667, -0.44598827, -0.47103143, -0.4984866, -0.5280283, -0.559114, -0.59120065, -0.62376297, -0.65642166, -0.68887436, -0.7208185, -0.7519693, -0.78221214, -0.8115235, -0.839879, -0.8672234, -0.8932216, -0.9173877, -0.9392363, -0.9582789, -0.9739766, -0.98576504, -0.9930836, -0.99543446, -0.99288875, -0.9858408, -0.9746934, -0.959853, -0.94171184, -0.9206539, -0.8970656, -0.87132764, -0.8437381, -0.81454027, -0.7839671, -0.75221866, -0.71925414, -0.68489045, -0.6489388, -0.6112349, -0.57191294, -0.5312845, -0.4896597, -0.447394, -0.40535906, -0.36473158, -0.32668006, -0.29230592, -0.2620922, -0.23614524, -0.21456765, -0.19745085, -0.1847412, -0.17629682, -0.17197888, -0.17164634, -0.17509009, -0.18294042, -0.19350097, -0.2070421, -0.2230696, -0.24098136, -0.26017603, -0.28005707, -0.30006287, -0.3196489, -0.33827037, -0.35541382, -0.3708345, -0.3844237, -0.39607406, -0.40569654, -0.41335812, -0.41920575, -0.42338738, -0.42605892, -0.42744604, -0.42781034, -0.4274132, -0.42651337, -0.42534998, -0.4241515, -0.42314544, -0.4225664, -0.4227188, -0.42394325, -0.4265831, -0.43096367, -0.43726695, -0.4455972, -0.45605907, -0.46874025, -0.48354506, -0.50028056, -0.5187521, -0.5387679, -0.5601599, -0.58277357, -0.6064534, -0.6310387, -0.65632135, -0.6820651, -0.708032, -0.7339808, -0.7596566, -0.78479624, -0.8091346, -0.83241946, -0.85454154, -0.86515886, -0.8854918, -0.90460426, -0.92252266, -0.9393819, -0.95533216, -0.97052455, -0.98512113, -0.9993086, -1.013277, -1.0272168, -1.0412219, -1.0551641, -1.0688841, -1.0822225, -1.0950212, -1.1071277, -1.1183891, -1.1286545, -1.1378762, -1.1462536, -1.1540223, -1.1614181, -1.1686246, -1.1757017, -1.1826912, -1.1896346, -1.1966047, -1.2037488, -1.2112249, -1.21919, -1.2278376, -1.2374535, -1.2483368, -999.0, -999.0, -1.2909749, -1.3086429, -1.3279532, -1.3487867, -1.3708576, -1.3938541, -1.4174656, -1.4413604, -1.4651519, -1.4884458, -1.5108485, -1.5320356, -1.5518636, -1.570219, -1.5885749, -1.6035513, -1.6170253, -1.6291449, -1.6400542, -1.6499614, -1.6592042, -1.6681353, -1.6771039, -1.6864386, -1.6964275, -1.707353, -1.7194974, -1.733064, -999.0, -999.0, -1.7825685, -1.8020582, -1.8230577, -1.8455708, -1.8696018, -1.8952842, -1.923037, -1.9533186, -1.9865881, -2.023254, -2.0636172, -2.107965, -2.156586, -2.2097278, -2.2675452, -2.330183, -2.3977904, -2.4705229, -2.5485442, -2.6320255, -2.721148, -2.8160539, -2.9167833, -3.0233717, -3.1358654, -3.2542558, -3.37838, -999.0, -3.643115, -3.7832398, -3.9277852, -4.076037, -999.0, -999.0, -4.5355964, -4.6911435, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -5.7271857, -5.8568487, -5.9789076, -6.092485, -6.1971765, -6.2926683, -6.3786654, -6.4550805, -6.5223346, -6.5809493, -6.631465, -6.6745105, -6.7109203, -6.741569, -6.7673364, -6.7891498, -6.808059, -6.8251343, -6.84144, -6.8579793, -6.875587, -6.8950686, -999.0, -999.0, -999.0, -7.004171, -7.040345, -7.08014, -7.1231585, -7.168941, -7.2170277, -7.2669287, -7.318065, -7.369842, -7.4216614, -7.4729033, -7.522896, -7.5709553, -7.6163974, -7.658585, -7.69702, -7.7312317, -7.7607546, -7.7851315, -7.8054795, -7.8176346, -7.823321, -7.8223567, -7.81507, -7.8018646, -999.0, -7.759501, -7.7318845, -7.701305, -7.668749, -7.635156, -999.0, -999.0, -7.536625, -7.5071154, -7.4800754, -7.4557867, -7.434523, -7.416654, -7.4027767, -7.3935137, -7.3894773, -7.391147, -7.3986883, -7.4122224, -7.4318757, -7.457717, -999.0, -999.0, -7.5714126, -7.6209645, -7.675814, -7.735506, -7.7995954, -7.867624, -7.9390836, -8.013462, -8.090246, -8.168831, -8.248371, -8.288221, -8.36751, -8.445514, -8.521766, -999.0, -999.0, -999.0, -8.80592, -8.871336, -8.934589, -8.995738, -9.054752, -9.111535, -9.165981, -999.0, -999.0, -9.314439, -9.358845, -9.400652, -9.43976, -9.476028, -9.509309, -9.539467, -9.566501, -9.590511, -9.611615, -9.6299515, -9.645885, -9.659955, -9.672704, -9.684688, -999.0, -9.708793, -9.722184, -9.737307, -9.75477, -9.775168, -9.799093, -999.0, -9.859319, -9.895517, -9.935469, -9.978934, -10.025506, -10.074644, -10.125802, -10.178456, -10.232374, -10.287562, -10.344037, -10.401822, -10.461008, -10.521747, -10.58419, -10.6484995, -10.714858, -10.783473, -10.854552, -10.928301, -11.004808, -11.084064, -11.166053, -11.250749, -999.0, -999.0, -999.0, -11.610499, -11.703373, -11.795952, -11.887309, -11.976498, -12.062653, -12.152981, -12.230199, -12.30195, -12.367734, -12.427249, -12.480209, -12.526364, -12.565752, -12.598616, -12.625218, -12.645845, -12.660948, -12.67109, -12.676842, -12.678772, -12.677429, -12.673348, -12.667057, -12.65907, -12.649799, -12.639585, -12.634226, -12.62321, -12.612013, -12.600754, -12.589523, -12.578412, -12.567508, -12.556909, -12.546709, -12.537004, -12.52792, -12.519686, -12.512542, -12.506728, -12.502445, -12.49979, -12.498844, -12.499682, -12.502352, -12.506812, -12.513007, -12.520882, -12.530369, -12.541362, -12.553748, -12.56742, -12.582224, -12.5978775, -12.614076, -12.630513, -12.646856, -12.662658, -12.677453, -12.690783, -12.702174, -12.711114, -12.717083, -12.719569, -12.718179, -12.7129, -12.703795, -12.690929, -12.674473, -12.654941, -12.6329155, -12.608972, -999.0, -999.0, -999.0, -12.498892, -12.467796, -12.435121, -12.4007225, -12.364466, -12.326299, -12.286464, -12.245262, -12.202987, -12.159946, -12.116516, -12.073081, -12.030013, -11.9876585, -11.946277, -11.906104, -11.86737, -11.830169, -11.794104, -11.758677, -11.723396, -11.687808, -11.651567, -11.614356, -11.575864, -11.535917, -11.49485, -11.453106, -11.411126, -11.36941, -11.328713, -11.289848, -11.2536125, -11.23344, -11.202675, -11.175659, -11.152603, -11.133694, -11.118756, -11.107347, -11.099021, -11.093334, -11.089737, -11.0876, -11.0863, -11.0852375, -999.0, -999.0, -999.0, -11.078286, -11.075164, -11.071315, -11.066679, -11.061199, -11.054836, -11.047572, -11.039385, -11.0302515, -11.020156, -11.009089, -10.997045, -10.984023, -10.970239, -10.956071, -10.941901, -10.928107, -10.915087, -10.9032545, -10.893021, -10.884783, -10.878748, -10.874964, -10.873475, -10.874321, -10.877401, -10.882494, -10.889379, -10.897832, -10.907594, -10.918369, -10.929863, -10.941785, -10.953923, -10.966132, -10.9782715, -10.990207, -11.001923, -11.013514, -11.025076, -11.036712, -11.048564, -11.060817, -11.073659, -11.08727, -11.101724, -11.116994, -11.133049, -11.149853, -11.167245, -11.184948, -11.202679, -11.220152, -11.236985, -11.252709, -11.266851, -11.27895, -11.28875, -11.296195, -11.301239, -11.303842, -11.30409, -11.302197, -11.298381, -11.292852, -11.285827, -11.28182, -11.272952, -11.263123, -11.252548, -11.241477, -11.230167, -11.218874, -11.207849, -11.197344, -11.187607, -11.178084, -11.170762, -11.164908, -11.160701, -11.158321, -11.157923, -11.159572, -11.163319, -11.169213, -11.177296, -11.187566, -11.200015, -11.214635, -11.231438, -11.250494, -11.271886, -11.295697, -11.322041, -11.351133, -11.383215, -11.418525, -11.457323, -11.499949, -11.54676, -11.598114, -11.654368, -11.715869, -11.782964, -11.856006, -11.935324, -12.021141, -12.113666, -12.213109, -12.319544, -12.4325285, -12.551505, -999.0, -12.80505, -12.937768, -13.072788, -13.2088175, -13.34458, -13.478899, -13.610612, -13.738542, -13.861549, -13.978681, -14.089022, -14.191649, -14.285784, -14.3712, -14.410612, -14.482792, -14.546067, -14.600707, -14.647306, -14.68648, -14.71885, -14.745003, -14.765485, -14.780846, -14.791631, -14.79819, -14.800688, -14.799276, -14.79411, -14.785262, -14.77273, -14.756507, -14.736585, -14.712937, -14.685521, -14.654288, -14.619198, -14.580359, -14.538037, -14.492498, -14.4440155, -14.39314, -14.340711, -14.287569, -14.234547, -14.182447, -14.132051, -14.084131, -14.039449, -13.998617, -13.962096, -13.930338, -13.903792, -13.882764, -13.867398, -13.8578415, -13.855286, -13.854658, -13.85982, -13.870521, -13.88651, -13.907513, -13.933133, -13.96294, -13.996505, -14.0334015, -14.077355, -14.119944, -14.164625, -14.2110405, -14.258965, -14.308205, -14.358566, -14.409882, -14.462073, -14.515087, -14.568869, -14.623382, -14.678664, -14.734771, -14.791756, -14.849676, -14.908593, -14.968573, -15.029676, -15.091953, -15.155379, -15.219916, -15.285527, -15.35217, -15.419801, -15.488372, -15.5578375, -15.628142, -15.699203, -15.7709255, -15.843218, -15.915996, -15.989195, -16.062761, -16.136637, -16.210764, -16.285065, -16.359453, -16.433846, -16.508114, -16.58194, -16.654953, -16.726788, -16.797085, -16.86555, -16.931894, -16.995832, -17.057123, -17.115707, -17.171572, -17.224707, -17.275146, -17.323124, -17.368923, -17.41283, -17.455143, -17.49621, -17.536396, -17.576065, -17.615553, -17.655062, -17.69476, -17.734814, -17.775358, -17.816399, -17.8579, -17.89983, -17.942156, -17.98486, -18.027924, -18.071335, -18.115068, -18.15905, -18.2032, -18.247429, -18.291653, -18.335781, -18.379725, -18.42339, -18.466696, -18.5096, -18.552076, -18.594093, -18.635628, -18.67665, -18.717134, -18.75706, -18.796394, -18.835098, -18.873129, -18.910439, -18.946997, -18.965, -19.000477, -19.035286, -19.069468, -19.103085, -19.136234, -19.169014, -19.20152, -19.233818, -19.265932, -19.301077, -19.332888, -19.364605, -19.396269, -19.427927, -19.459625, -19.491398, -19.523272, -19.555277, -19.587435, -19.61975, -19.652191, -19.684732, -19.717352, -19.75008, -19.783016, -19.816256, -19.849897, -19.884012, -19.918646, -19.953844, -19.98965, -20.026085, -20.063139, -20.100811, -20.139091, -20.177986, -20.217508, -20.257675, -20.298502, -20.339998, -20.382174, -20.42503, -20.468578, -20.512825, -20.557777, -20.603449, -20.649845, -20.696957, -20.74475, -20.793188, -20.84224, -20.891815, -20.941776, -20.991982, -21.042286, -21.092566, -21.142717, -21.19264, -21.24223, -21.29137, -21.339937, -21.387802, -21.434834, -21.480883, -21.525776, -21.569338, -21.611385, -21.651512, -21.689035, -21.723257, -21.753496, -21.779661, -21.802383, -21.82233, -21.840172, -21.856573, -21.87219, -21.88768, -21.903692, -21.920704, -21.93898, -21.948671, -21.96931, -21.991823, -22.016354, -22.043026, -22.071957, -22.103247, -22.136873, -22.172773, -22.210882, -22.251133, -22.29342, -22.337627, -22.383638, -22.431335, -22.480595, -22.531284, -22.58328, -22.63645, -22.690634, -22.74566, -22.801365, -22.857578, -22.91415, -22.97093, -23.027775, -23.084543, -23.141132, -23.197456, -23.253426, -23.308949, -23.36389, -23.418108, -23.471457, -23.5238, -23.575048, -23.625135, -23.673992, -23.721565, -23.767889, -23.813028, -23.861397, -23.904268, -23.946144, -23.987068, -24.027082, -24.066233, -24.104574, -24.142157, -24.179037, -24.215271, -24.250938, -24.286121, -24.320902, -24.355364, -24.3896, -24.423708, -24.457779, -24.491903, -24.526133, -24.560513, -24.595083, -24.629887, -24.664927, -24.7002, -24.735703, -24.771431, -24.807367, -24.843487, -24.87977, -24.916193, -24.952719, -24.989305, -25.025915, -25.062513, -25.099113, -25.135736, -25.17241, -25.209167, -25.246107, -25.283352, -25.32102, -25.359226, -25.398048, -25.437561, -25.477829, -25.518919, -25.560848, -25.603628, -25.647264, -25.69176, -25.737091, -25.783228, -25.830137, -25.877785, -25.926123, -25.975094, -26.024645, -26.074726, -26.125334, -26.176474, -26.228151, -26.280373, -26.333103, -26.386301, -26.439922, -26.493923, -26.548256, -26.602879, -26.657745, -26.712797, -26.767897, -26.822876, -26.877563, -26.931772, -26.985188, -27.037443, -27.088173, -27.137012, -27.183592, -27.227547, -27.268509, -27.306145, -27.340317, -27.370974, -27.398062, -27.421583, -27.441883, -27.459438, -27.47473, -27.488247, -27.500525, -27.512112, -27.523558, -27.535412, -27.54819, -27.562407, -27.57857, -27.597158, -27.618467, -27.642714, -27.67011, -27.700846, -27.73849, -27.776093, -27.816818, -27.86054, -27.907015, -27.955952, -28.007065, -28.060057, -28.114586, -28.170298, -28.226837, -28.283848, -28.340973, -28.397852, -28.454126, -28.509453, -28.563557, -28.616188, -28.6671, -28.716068, -28.762974, -28.80774, -28.850292, -28.89058, -28.928705, -28.964828, -28.999102, -29.031702, -29.062902, -29.093016, -29.122349, -29.15121, -29.179876, -29.208614, -29.23769, -29.26737, -29.297916, -29.329594, -29.362661, -29.397354, -29.433754, -29.471878, -29.51175, -29.553362, -29.596586, -29.641233, -29.687117, -29.734058, -29.781933, -29.83063, -29.880037, -29.930037, -29.980427, -30.030973, -30.081444, -30.131607, -30.18122, -30.23004, -30.277826, -30.324354, -30.369524, -30.413294, -30.455618, -30.496471, -30.535963, -30.57426, -30.61153, -30.647943, -30.683704, -30.71903, -30.754139, -30.789248, -30.824547, -30.842327, -30.878258, -30.91484, -30.952164, -30.990173, -31.028795, -31.06796, -31.107595, -31.14762, -31.187954, -31.208212, -31.248865, -31.28969, -31.330675, -31.37182, -31.41311, -31.454475, -31.495817, -31.537039, -31.578035, -31.622654, -31.662558, -31.70161, -31.7396, -31.776264, -31.811335, -31.844543, -31.875635, -31.904455, -31.930883, -31.954802, -31.976126, -31.994968, -32.01152, -32.02597, -32.038536, -32.049576, -32.05952, -32.068787, -32.0778, -32.082344, -32.09175, -32.101936, -32.113316, -32.12628, -32.141216, -32.158493, -32.178486, -32.201496, -32.227703, -32.257275, -32.273373, -32.30826, -32.34655, -32.38796, -32.4322, -32.478973, -32.527824, -32.578255, -32.62976, -32.681835, -32.733932, -32.75982, -32.81091, -32.86064, -32.90852, -32.95417, -32.997215, -33.037285, -33.07411, -33.107563, -33.13753, -33.163902, -33.18661, -33.205647, -33.221012, -33.232704, -33.24055, -33.244125, -33.242973, -33.236645, -33.22527, -33.209892, -33.191658, -33.171696, -33.15117, -33.131256, -33.11315, -33.098022, -33.08663, -33.07902, -33.075165, -33.075035, -33.078465, -33.08505, -33.094357, -33.10596, -33.11941, -33.134216, -33.149895, -33.16595, -33.181946, -33.1975, -33.212246, -33.2192, -33.232063, -33.243385, -33.253033, -33.26087, -33.26678, -33.2707, -33.272606, -33.27248, -33.2703, -33.26844, -33.26319, -33.255913, -33.246624, -33.235382, -33.222355, -33.207703, -33.191605, -999.0, -999.0, -999.0, -999.0, -33.104115, -33.081856, -33.058823, -33.03515, -33.010952, -32.98629, -32.961178, -32.935627, -32.922695, -32.896523, -32.88062, -32.853786, -32.82654, -32.7989, -32.771008, -32.743042, -32.71519, -32.687653, -32.660667, -32.634518, -32.609467, -32.58577, -32.563488, -32.542625, -32.523167, -32.505104, -32.488358, -32.472824, -32.4584, -32.444984, -32.432495, -32.420856, -32.40999, -32.399803, -32.390133, -32.380768, -32.371506, -32.362125, -32.352375, -32.341984, -32.330677, -32.324593, -32.311466, -32.296986, -32.28107, -32.26364, -32.244686, -32.224342, -32.20274, -32.180027, -32.15641, -32.132225, -32.107822, -32.083546, -32.059757, -32.03685, -32.015224, -31.995272, -31.977304, -31.961494, -31.947998, -31.936966, -31.928417, -31.922113, -31.917797, -31.915203, -31.91396, -31.913494, -31.913206, -31.912504, -31.910898, -31.908102, -31.903856, -31.897896, -31.890076, -31.880466, -31.869162, -31.85626, -31.841896, -31.826284, -31.809654, -31.792229, -31.783287, -31.765083, -31.746634, -31.728155, -31.709856, -31.691883, -31.674347, -31.657358, -31.641018, -31.625324, -31.61022, -31.595646, -31.58154, -31.567787, -31.554247, -31.540777, -31.527235, -31.513447, -31.49923, -31.484398, -31.467175, -31.450651, -31.433334, -31.415257, -31.396456, -31.377016, -31.357042, -31.336637, -31.315908, -31.294937, -31.273808, -31.252596, -31.231384, -31.21024, -31.189228, -31.168415, -31.147863, -31.127588, -31.107595, -31.087881, -31.068453, -31.049345, -31.039927, -31.021389, -31.003292, -30.98567, -30.968542, -30.951916, -30.935806, -30.920221, -30.90516, -30.89062, -30.876595, -30.863073, -30.850008, -30.837353, -30.825058, -30.813038, -30.801136, -30.789186, -30.777021, -30.764547, -30.751787, -30.73878, -30.725563, -30.712208, -30.698835, -30.685577, -30.67256, -30.659899, -30.647669, -30.635944, -30.624802, -30.6143, -30.604473, -30.595352, -30.586967, -30.57936, -30.572596, -30.56674, -30.561863, -30.55803, -30.555313, -30.553783, -30.553486, -30.553865, -30.555553, -30.55855, -30.562849, -30.56844, -30.575233, -30.583101, -30.591908, -30.601496, -30.611412, -30.621048, -30.62979, -30.637045, -30.642427, -30.645668, -30.646494, -30.644701, -30.640717, -30.635326, -30.629326, -30.623476, -30.618202, -30.61374, -30.610323, -30.60817, -30.607355, -30.607874, -30.609718, -30.612879, -30.6173, -30.622904, -30.62961, -30.637339, -30.645952, -30.655287, -30.665176, -30.675457, -30.685966, -30.69761, -30.708101, -30.718342, -30.728163, -30.737389, -30.745846, -30.753366, -30.759825, -30.765114, -30.769129, -30.771765, -30.772924, -30.77292, -30.771687, -30.768736, -30.76419, -30.758568, -30.752432, -30.746347, -30.740978, -30.737188, -30.735865, -30.737888, -30.744019, -30.754765, -30.770613, -30.79204, -30.819054, -30.850727, -30.886028, -30.923922, -30.96355, -31.004412, -31.046041, -31.087976, -31.129847, -31.171474, -31.212698, -31.253363, -31.293373, -31.332758, -31.371565, -31.409842, -31.447638, -31.485014, -31.522028, -31.55874, -31.59522, -31.631554, -31.667822, -31.704113, -31.740513, -31.77711, -31.813986, -31.85123, -31.888931, -31.927189, -31.966105, -32.00578, -32.046303, -32.087746, -32.130165, -32.173634, -32.195766, -32.240784, -32.2867, -32.333397, -32.38076, -32.428665, -32.476986, -32.525604, -32.574394, -32.623276, -32.672188, -32.721066, -32.76985, -32.818474, -32.86685, -32.914913, -32.962585, -33.00986, -33.056767, -33.10334, -33.149605, -33.17261, -33.21834, -33.263626, -33.30839, -33.35257, -33.39607, -33.43879, -33.480648, -33.521564, -33.561504, -33.60044, -33.638336, -33.675186, -33.71102, -33.745884, -33.77981, -33.812866, -33.84513, -33.87671, -33.90769, -33.93816, -33.968174, -33.99778, -34.027027, -34.055943, -34.084488, -34.112625, -34.140312, -34.167503, -34.194168, -34.22286, -34.248325, -34.2732, -34.297546, -34.32143, -34.344917, -34.368073, -34.390965, -34.413654, -34.436203, -34.45866, -34.48103, -34.503315, -34.52552, -34.54764, -34.56967, -34.591606, -34.61343, -34.635136, -34.656677, -34.678013, -34.69911, -34.709553, -34.73026, -34.75074, -34.77103, -34.791164, -34.811184, -34.831135, -34.851063, -34.87102, -34.8911, -34.911434, -34.93214, -34.953346, -34.97515, -34.99764, -35.020897, -35.045, -35.069977, -35.095814, -35.122498, -35.15002, -35.17836, -35.2075, -35.237415, -999.0, -999.0, -35.331173, -35.363297, -35.395596, -35.427963, -35.46033, -35.492615, -35.508705, -35.54075, -35.57262, -999.0, -999.0, -999.0, -999.0, -999.0, -35.761524, -35.777355, -35.809273, -35.841663, -35.874695, -35.908535, -35.94326, -35.9789, -36.015484, -36.05303, -36.091522, -36.13094, -36.15098, -36.191715, -36.23331, -36.27583, -36.31935, -36.363953, -36.409653, -36.45632, -36.5038, -36.551926, -36.60051, -36.624874, -36.67355, -36.721874, -36.769516, -36.816032, -36.86092, -36.903652, -36.943745, -36.980965, -999.0, -37.049656, -37.07787, -37.10387, -37.128708, -37.15344, -37.179066, -37.2061, -37.23476, -37.265255, -37.29778, -37.332367, -37.350414, -37.387966, -37.42741, -37.46862, -37.511353, -37.555336, -37.600315, -37.646065, -37.692486, -37.739494, -37.787003, -37.81092, -37.85911, -37.90779, -37.957, -38.00678, -38.057144, -38.108105, -38.15968, -38.211872, -38.264713, -38.318237, -38.345264, -38.399868, -38.455227, -38.511345, -38.56822, -38.625847, -38.684246, -38.743492, -38.803665, -38.86484, -38.895832, -38.958645, -39.022606, -39.087757, -39.15414, -39.221718, -39.290413, -39.360146, -39.430824, -39.502262, -39.57421, -39.646423, -39.718624, -39.79029, -39.860706, -39.92917, -39.994984, -40.05784, -40.11768, -40.174458, -40.228153, -40.253925, -40.303688, -40.35155, -40.39809, -40.44376, -40.48863, -40.532707, -40.575996, -40.61851, -40.66027, -40.701294, -40.741604, -40.781208, -40.820076, -40.858166, -40.89545, -40.931892, -40.96751, -41.002316, -41.036327, -41.06958, -41.102165, -41.13419, -41.165752, -41.196964, -41.22795, -41.25884, -41.28976, -41.320854, -41.352306, -41.38431, -41.40058, -41.43377, -41.467915, -41.50307, -41.5393, -41.57665, -41.61508, -41.65449, -41.69477, -41.735798, -41.756542, -41.79837, -41.840473, -41.882637, -41.924664, -41.96635, -42.00751, -42.047947, -42.087486, -42.12602, -42.16713, -42.203243, -42.23807, -42.2716, -42.303802, -42.334663, -42.36418, -42.392384, -42.4193, -42.444965, -42.469433, -42.48126, -42.504158, -42.52618, -42.547443, -42.568066, -42.58815, -42.607796, -42.627094, -42.64608, -42.664722, -42.683, -42.691994, -42.709675, -42.726933, -42.743744, -42.76009, -42.775948, -42.79127, -42.806007, -42.820118, -42.833557, -42.846325, -42.852455, -42.86421, -42.87529, -42.8858, -42.895912, -42.905807, -42.91567, -42.925735, -42.936287, -42.947613, -42.95999, -42.96664, -42.980934, -42.996662, -43.013947, -43.03287, -43.053394, -43.075447, -43.09896, -43.12388, -43.150166, -43.177795, -43.1921, -43.221687, -43.252563, -43.28472, -43.318172, -43.35291, -43.388943, -43.42627, -43.464897, -43.504826, -43.54603, -43.588444, -43.63202, -43.676693, -43.72235, -43.76883, -43.81597, -43.863617, -43.91158, -43.95967, -44.007698, -44.05546, -44.102753, -44.149353, -44.19504, -44.239594, -44.282803, -44.324474, -44.364414, -44.402435, -44.43847, -44.45575, -44.488865, -44.520084, -44.54948, -44.577232, -44.603542, -44.628616, -44.65266, -44.67587, -44.700665, -44.722744, -44.744583, -44.76635, -44.788216, -44.810352, -44.832897, -44.855892, -44.879368, -44.90335, -44.92785, -44.94027, -44.96541, -44.990883, -45.016617, -45.04257, -45.068718, -45.095043, -45.12153, -45.148193, -45.175095, -45.202282, -45.22981, -45.25772, -45.28605, -45.314827, -45.34409, -45.37381, -45.403946, -45.434437, -45.46523, -45.49625, -45.511818, -45.543015, -45.57421, -45.605343, -45.63638, -45.667305, -45.698112, -45.72876, -45.759136, -45.789116, -45.803917, -45.83307, -45.861576, -45.889427, -45.916615, -45.94312, -45.968983, -45.99427, -46.01904, -46.04336, -46.067314, -46.09098, -46.102734, -999.0, -46.149452, -46.172764, -46.19613, -46.219612, -46.243267, -46.26709, -46.29108, -46.31523, -46.33953, -46.363976, -46.388557, -46.413273, -46.43812, -46.463135, -46.488342, -46.51378, -46.53947, -46.56541, -46.57847, -46.60475, -46.63124, -46.657936, -46.684834, -46.711937, -46.739246, -46.766777, -46.794544, -46.82257, -999.0, -46.879436, -46.893795, -46.922634, -46.951588, -46.980618, -47.009735, -47.038975, -47.068367, -47.097935, -47.12766, -47.157513, -47.187477, -47.21752, -47.247623, -999.0, -999.0, -999.0, -999.0, -47.398388, -47.42872, -47.4592, -47.477577, -47.508373, -47.539406, -47.5707, -47.602314, -47.63432, -47.66678, -47.69977, -47.73338, -47.767693, -47.78514, -47.820686, -47.857143, -47.89451, -47.93276, -47.97187, -48.011818, -48.052517, -48.0939, -48.13588, -48.178387, -48.221413, -48.26494, -48.308952, -48.35344, -999.0, -999.0, -999.0, -999.0, -999.0, -48.626335, -48.649223, -48.69492, -48.740368, -999.0, -999.0, -999.0, -48.915794, -48.957066, -999.0, -999.0, -49.071533, -49.10609, -49.138687, -49.16923, -49.197525, -49.223278, -49.246204, -49.266033, -999.0, -49.29728, -49.30972, -49.320717, -49.330692, -49.33998, -49.348915, -49.35782, -49.36687, -49.37611, -49.385582, -49.39531, -49.40529, -49.415443, -49.425713, -49.430866, -49.441185, -49.451515, -49.46185, -49.472187}
rh =
  {47.3, 45.565132, 45.47368, 45.383923, 45.296703, 45.212746, 45.132256, 45.055317, 44.982002, 44.912464, 44.847137, 44.786533, 44.731167, 44.68159, 44.63854, 44.602783, 44.575108, 44.556248, 44.54678, 44.547226, 44.558117, 44.579967, 44.613274, 44.658504, 44.71615, 44.78668, 44.870564, 44.96827, 45.08026, 45.206894, 45.348026, 45.50338, 45.67267, 45.855442, 46.05048, 46.256332, 46.471558, 46.69455, 46.922943, 47.15416, 47.385624, 47.614708, 47.83853, 48.054157, 48.258644, 48.449394, 48.62546, 48.7864, 48.931763, 49.061035, 49.173374, 49.26785, 49.34352, 49.399334, 49.433628, 49.44455, -999.0, 49.389168, 49.321125, 49.226383, 49.09165, 48.941406, 48.76357, 48.55672, 48.31944, 48.0505, 47.749462, 47.416065, 47.05005, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 40.820965, -999.0, -999.0, -999.0, 38.43226, 37.850838, 37.28152, 36.72659, 36.188313, 35.668633, 35.1681, 34.68688, 34.225155, 33.78318, 33.361553, 32.960976, 32.582138, 32.225437, 31.889942, 31.574358, 31.277395, 30.99771, 30.733713, 30.483753, -999.0, 30.019575, 29.803572, 29.598104, 29.403107, 29.21851, 29.044245, 28.880243, 28.726435, 28.582766, -999.0, -999.0, 28.212725, 28.109787, 28.017084, 27.934635, 27.862455, 27.800465, 27.748137, 27.70481, 27.669819, 27.642431, 27.621561, 27.606018, 27.59461, 27.586231, 27.580206, 27.575993, 27.573048, 27.570992, 27.570246, 27.571493, 27.575415, 27.582653, 27.593678, 27.6089, 27.628733, 27.653475, 27.682858, 27.716425, 27.753714, 27.794195, 27.836918, 27.880806, 27.924774, 27.967735, 28.008574, 28.046156, 28.079353, 28.107298, 28.130558, 28.150194, 28.167269, 28.182804, 28.197617, 28.21397, 28.2297, 28.247011, 28.266588, 28.289106, 28.315239, 28.345598, 28.380535, 28.42033, 28.465265, 28.515427, 28.570055, 28.628159, 28.68875, 28.750795, 28.813084, 28.874353, 28.933344, 28.988924, 29.040575, 29.087944, 29.130674, 29.168499, 29.201529, 29.229982, 29.254082, 29.273985, 29.28958, 29.300673, 29.307072, 29.308832, 29.307175, 29.303658, 29.299847, 29.297272, 29.29731, 29.301292, 29.310555, 29.326159, 29.347878, 29.375084, 29.407152, 29.443161, 29.48073, 29.517025, 29.549213, 29.574688, 29.591995, 29.600039, 29.597725, 29.584269, 29.560484, 29.527683, 29.487188, 29.440264, 29.387915, 29.33106, 29.270618, 29.207413, 29.14177, 29.073847, 29.003807, 28.931805, 28.85798, 28.782463, 28.705387, 28.626902, 28.547277, 28.466825, 28.38585, 28.30471, 28.22399, 28.144356, 28.066483, 27.990847, 27.916845, 27.8435, 27.769829, 27.694862, 27.617691, 27.537424, 27.453175, 27.364296, 27.271545, 27.176193, 27.079508, 26.982855, 26.88817, 26.797594, 26.713268, 26.637157, 26.570139, 26.512686, 26.465271, 26.42825, 26.401253, 26.383642, 26.374775, 26.374071, 26.381332, 26.396511, 26.41956, 26.450611, 26.490967, 26.548208, 26.613832, 26.694208, 26.791046, 26.906048, 27.040913, 27.197187, 27.37567, 27.57693, 27.80154, 28.049911, 28.321655, 28.616146, 28.932753, 29.27067, 29.628212, 30.003416, 30.394327, -999.0, -999.0, 31.641077, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 35.94199, -999.0, -999.0, 37.05139, -999.0, -999.0, -999.0, -999.0, -999.0, 38.84007, 39.080685, -999.0, -999.0, -999.0, -999.0, -999.0, 40.14225, -999.0, -999.0, -999.0, -999.0, 40.4452, 40.436073, 40.402924, 40.34553, 40.2643, 40.159843, 40.032772, 39.883865, 39.7149, 39.528008, 39.325325, 39.109173, 38.882954, 38.650482, 38.415585, 38.18186, 37.95163, 37.72672, 37.50895, 37.299942, 37.100044, 36.90911, -999.0, -999.0, 36.386253, 36.223362, 36.062233, 35.900497, 35.736183, 35.56745, 35.39248, 35.209675, 35.019012, 34.82111, 34.616585, 34.406197, 34.1917, 33.975246, 33.75899, 33.54501, 33.334873, 33.129917, 32.931488, 32.740856, -999.0, -999.0, -999.0, 32.0694, 31.928284, 31.801132, 31.68998, 31.588478, 31.516357, 31.464342, 31.433308, 31.42381, 31.434677, 31.464155, 31.51049, 31.571903, 31.646448, 31.732124, 31.826935, -999.0, -999.0, 32.14495, 32.25456, 32.362183, 32.465828, -999.0, -999.0, -999.0, -999.0, 32.863266, 32.910908, 32.946712, 32.97162, 32.987, 32.994247, 32.994785, 32.990295, 32.98255, 32.97332, 32.964237, 32.956123, 32.94947, 32.94479, 32.9426, 32.943516, 32.948185, 32.95726, 32.97141, 32.99135, 33.017834, 33.051613, 33.093426, 33.143963, 33.203888, 33.273872, 33.354553, 33.446396, 33.549793, 33.66514, 33.792778, 33.932762, 34.08502, 34.249466, 34.425922, 34.613426, 34.810703, 35.016476, 35.229515, 35.448902, 35.67384, 35.903534, 36.13716, 36.373695, 36.612026, 36.851032, 37.089645, 37.327038, 37.56249, 37.79529, 38.024826, 38.251213, 38.474888, 38.69629, 38.915897, 39.134514, 39.353085, 39.57256, 39.793957, 40.018887, 40.2492, 40.48676, 40.73322, 40.988636, 41.252365, 41.52374, 41.802044, 42.086124, 42.374615, 42.666157, -999.0, -999.0, 43.57786, 43.872364, 44.16616, 44.458878, 44.750206, 45.039825, 45.32721, 45.610573, 45.887676, 46.15628, 46.41447, 46.66227, 46.90042, 47.129677, 47.350845, 47.565136, 47.773914, 47.978535, 48.18036, 48.38075, 48.58106, 48.782654, 48.986786, 49.194065, 49.404858, 49.619522, 49.83834, 50.061058, 50.28722, 50.516365, 50.74785, 50.979805, -999.0, -999.0, 51.655113, 51.86632, 52.067924, 52.25849, 52.43677, 52.602795, 52.757103, 52.900246, 53.032852, 53.156044, 53.27116, 53.379528, 53.482544, 53.581993, 53.67983, 53.778004, 53.878395, 53.982327, 54.09088, 54.20515, 54.326088, 54.453766, 54.587852, 54.728024, 54.873947, 55.02528, 55.18167, 55.342766, 55.50815, 55.67682, 55.84754, 56.019073, 56.19023, 56.360332, 56.528908, 56.6955, 56.85969, 57.021416, 57.180786, 57.3379, 57.492657, 57.64335, 57.7875, 57.922634, 58.04615, 58.15447, 58.243538, 58.309303, 58.347782, 58.35557, 58.329563, 58.266647, -999.0, -999.0, 57.835667, 57.609776, -999.0, -999.0, -999.0, -999.0, -999.0, 55.447544, 54.972534, -999.0, -999.0, 53.40872, 52.856216, 52.297245, -999.0, -999.0, 50.64051, -999.0, 49.616924, 49.146824, 48.7098, 48.30959, 47.91605, 47.60256, 47.332054, 47.10532, 46.92281, 46.782707, 46.682255, 46.618683, 46.589203, 46.590775, 46.620277, 46.674576, 46.750607, 46.845802, 46.957798, 47.084225, 47.22274, 47.371048, 47.5269, 47.688038, 47.852314, 48.01835, 48.185097, 48.351524, 48.51685, 48.682198, 48.849564, 49.020927, 49.198303, 49.38386, 49.57984, 49.788483, 50.01184, 50.25055, 50.50458, 50.773903, 51.0582, 51.35485, 51.660168, 51.970455, 52.28206, 52.591606, 52.89587, 53.19162, 53.47582, 53.7469, -999.0, -999.0, -999.0, 54.68373, 54.877693, 55.054565, 55.214134, 55.358265, 55.48987, 55.61186, 55.727062, 55.837616, 55.945293, 56.05186, 56.158905, 56.266373, 56.37336, 56.47897, -999.0, -999.0, 56.781715, 56.87773, 56.97142, 57.063564, 57.15529, 57.247734, 57.341915, 57.43774, 57.53453, 57.631596, 57.728165, 57.822643, 57.912994, -999.0, 58.073326, 58.141506, 58.202797, 58.25828, 58.309093, 58.35661, 58.40237, 58.44791, 58.49477, 58.544422, 58.598328, 58.65794, 58.73172, 58.806828, 58.88968, 58.98037, 59.07881, 59.18364, 59.29292, 59.4047, 59.517193, 59.629597, 59.741573, 59.8528, 59.963013, 60.072582, 60.182156, 60.292374, 60.40388, 60.51727, 60.633114, 60.751984, 60.874496, 61.00157, 61.134285, 61.273712, 61.420826, 61.57581, 61.73847, 61.908596, 62.08586, 62.268833, 62.455547, 62.64404, 62.83242, 63.019444, 63.20417, 63.38567, 63.563057, 63.73589, 63.903934, 64.06696, 64.224815, 64.37794, 64.52706, 64.67295, 64.81627, 64.95703, 65.09491, 65.22958, 65.36081, 65.48914, 65.61555, 65.741005, 65.8664, 65.991844, 66.11702, 66.241615, 66.36528, 66.48731, 66.6068, 66.72285, 66.83471, 66.943184, 67.0499, 67.1565, 67.26471, 67.37692, 67.49593, 67.62455, 67.76547, 67.9206, 68.091385, 68.27925, 68.48556, 68.71071, 68.954575, 69.21704, 69.49781, 69.79485, 70.10515, 70.42565, 70.75345, 71.08684, 71.42483, 71.76646, 72.110725, 72.45656, 72.8028, 73.14832, 73.49177, 73.82975, 74.157616, 74.470695, 74.76453, 75.03687, 75.286865, 75.51368, 75.71653, 75.89537, 76.05061, 76.18267, 76.29199, 76.379234, 76.45069, 76.49426, 76.518524, 76.52613, 76.52056, 76.505295, 76.48377, 76.4591, 76.43422, 76.41207, 76.39543, 76.38555, 76.38294, 76.3881, 76.40146, 76.42286, 76.45185, 76.487976, 76.530716, 76.579056, 76.63169, 76.68732, 76.74463, 76.80221, 76.858574, 76.91226, 76.961754, 77.00521, 77.04062, 77.065956, 77.07931, 77.07961, 77.066284, 77.03873, 76.9965, 76.94027, 76.87136, 76.791115, 76.70083, 76.6018, 76.49527, 76.38249, 76.26475, 76.14362, 76.02091, 75.89837, 75.777794, 75.661026, 75.54996, 75.44648, 75.35238, 75.26824, 75.22987, 75.16049, 75.10081, 75.05043, 75.008316, 74.97333, 74.94434, 74.920235, 74.89989, 74.882195, 74.86606, 74.850945, 74.837654, 74.82718, 74.82051, 74.818695, 74.822914, 74.83436, 74.85422, 74.8831, 74.92025, 74.96469, 75.01545, 75.07183, 75.13377, 75.201324, 75.27451, 75.35305, 75.435844, 75.521675, 75.609314, 75.69741, 75.784225, 75.868, -999.0, -999.0, 76.08638, 76.14687, 76.20133, 76.2502, 76.294716, 76.336296, 76.37633, 76.41632, 76.45809, 76.50347, 76.55433, 76.61208, 76.67707, 76.749435, 76.83772, 76.92552, 77.01909, 77.11689, 77.2174, 77.31869, 77.418015, 77.51254, 77.59941, 77.67589, 77.73947, 77.787674, 77.818016, 77.828896, -999.0, -999.0, 77.74798, 77.685265, 77.607445, 77.51685, 77.41582, 77.30587, 77.18684, 77.05828, 76.9198, 76.77087, 76.61073, 76.43863, 76.25377, 76.0552, 75.84156, 75.61141, 75.363335, 75.09578, 74.806885, 74.49477, 74.15752, 73.79346, 73.40139, 72.98017, 72.52867, 72.04635, 71.534, -999.0, 70.42323, 69.82774, 69.21021, 68.57503, -999.0, -999.0, 66.60958, 65.95214, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 61.853256, 61.39222, 60.973465, 60.59951, 60.27048, 59.98612, 59.746162, 59.549633, 59.393696, 59.275223, 59.191074, 59.13791, 59.111847, 59.108906, 59.12511, 59.156414, 59.19854, 59.24719, 59.298058, 59.3471, 59.39097, 59.42644, -999.0, -999.0, -999.0, 59.435043, 59.39994, 59.350006, 59.28714, 59.21352, 59.131313, 59.042862, 58.95098, 58.85856, 58.76849, 58.683662, 58.606922, 58.54112, 58.4891, 58.453457, 58.436043, 58.438576, 58.46277, 58.51049, 58.592888, 58.697563, 58.833035, 59.000626, 59.199272, 59.42757, -999.0, 59.96666, 60.270916, 60.592335, 60.926365, 61.26869, -999.0, -999.0, 62.30797, 62.646706, 62.977455, 63.298466, 63.60798, 63.90359, 64.181335, 64.437, 64.66639, 64.86578, 65.03264, 65.16462, 65.25935, 65.31498, -999.0, -999.0, 65.24111, 65.135216, 64.99043, 64.80876, 64.59221, 64.34295, 64.063515, 63.756523, 63.424583, 63.070805, 62.69958, 62.508873, 62.120132, 61.725365, 61.327564, -999.0, -999.0, -999.0, 59.744225, 59.358135, 58.978096, 58.6051, 58.24054, 57.886097, 57.543457, -999.0, -999.0, 56.603817, 56.326263, 56.069702, 55.836105, 55.62751, 55.44594, 55.293327, 55.170162, 55.07586, 55.0098, 54.97128, 54.958183, 54.967346, 54.995575, 55.03965, -999.0, 55.16085, 55.23034, 55.300655, 55.36807, 55.428917, 55.47953, -999.0, 55.537693, 55.54324, 55.532772, 55.5061, 55.46387, 55.407402, 55.338036, 55.257046, 55.16475, 55.06068, 54.94435, 54.815273, 54.67302, 54.517193, 54.347404, 54.16328, 53.96465, 53.7515, 53.523846, 53.281708, 53.025517, 52.756058, 52.47411, 52.18052, -999.0, -999.0, -999.0, 50.933235, 50.617313, 50.307632, 50.00884, 49.72553, 49.46155, 49.197304, 48.984264, 48.80027, 48.647038, 48.525333, 48.435925, 48.379475, 48.35544, 48.362434, 48.399055, 48.46385, 48.55473, 48.669155, 48.804585, 48.958477, 49.128487, 49.312393, 49.507984, 49.713074, 49.925934, 50.145153, 50.256714, 50.48286, 50.71209, 50.94378, 51.177425, 51.41252, 51.648552, 51.884983, 52.121284, 52.356922, 52.591206, 52.823017, 53.05114, 53.27436, 53.491585, 53.702023, 53.90495, 54.09964, 54.28552, 54.46247, 54.630463, 54.789463, 54.93955, 55.08115, 55.21476, 55.340878, 55.460224, 55.57426, 55.684586, 55.79281, 55.90066, 56.010345, 56.124134, 56.244316, 56.373154, 56.512863, 56.665657, 56.833744, 57.018814, 57.220837, 57.439445, 57.67426, 57.924507, 58.188076, 58.46259, 58.745655, -999.0, -999.0, -999.0, 59.947784, 60.26794, 60.597263, 60.93658, 61.28672, 61.64808, 62.01955, 62.39968, 62.787037, 63.18008, 63.576958, 63.975742, 64.374504, 64.77141, 65.164925, 65.55361, 65.93601, 66.311356, 66.68136, 67.048294, 67.41446, 67.782005, 68.15258, 68.52773, 68.90899, 69.29727, 69.69122, 70.08891, 70.48841, 70.88752, 71.28292, 71.67104, 72.04832, 72.26809, 72.62235, 72.96085, 73.282745, 73.587296, 73.875534, 74.1498, 74.41249, 74.66604, 74.913536, 75.15861, 75.40489, 75.65591, -999.0, -999.0, -999.0, 76.727005, 77.01206, 77.30295, 77.59871, 77.89844, 78.201294, 78.50657, 78.81354, 79.12149, 79.43016, 79.73962, 80.04993, 80.3611, 80.671776, 80.97947, 81.281654, 81.57581, 81.8593, 82.129364, 82.383255, 82.6183, 82.83328, 83.02818, 83.20303, 83.357925, 83.49359, 83.61139, 83.71268, 83.79882, 83.87121, 83.93125, 83.980354, 84.01992, 84.05127, 84.07562, 84.09421, 84.10823, 84.11857, 84.12578, 84.13043, 84.13307, 84.13442, 84.13532, 84.13661, 84.139145, 84.143906, 84.151985, 84.16448, 84.18251, 84.20705, 84.239, 84.27926, 84.32876, 84.38898, 84.46195, 84.54975, 84.65436, 84.77653, 84.91574, 85.07146, 85.24308, 85.42903, 85.62676, 85.83368, 86.0472, 86.26493, 86.37469, 86.59459, 86.8132, 87.02844, 87.2388, 87.44291, 87.63939, 87.82705, 88.00548, 88.174484, 88.34926, 88.49798, 88.637535, 88.76858, 88.89172, 89.007645, 89.1171, 89.22087, 89.319725, 89.41436, 89.50517, 89.59251, 89.67671, 89.757835, 89.83503, 89.907234, 89.97339, 90.03219, 90.0815, 90.118965, 90.14229, 90.14901, 90.136314, 90.101295, 90.04104, 89.95275, 89.83409, 89.68279, 89.49658, 89.273605, 89.013435, 88.71594, 88.381004, 88.00922, 87.60372, 87.16821, -999.0, 86.222496, 85.72253, 85.212906, 84.70009, 84.1903, 83.689, 83.201485, 82.73305, 82.28881, 81.87326, 81.49074, 81.145584, 80.84153, 80.57999, 80.46543, 80.26927, 80.117714, 80.010056, 79.94414, 79.91774, 79.92864, 79.97455, 80.05307, 80.16183, 80.298454, 80.46122, 80.64901, 80.86073, 81.095314, 81.35182, 81.62946, 81.92747, 82.24503, 82.5814, 82.935776, 83.30738, 83.6954, 84.098434, 84.514465, 84.94143, 85.37724, 85.81863, 86.2611, 86.7001, 87.13109, 87.54986, 87.95255, 88.33535, 88.69445, 89.02709, 89.33163, 89.60647, 89.850044, 90.06168, 90.241684, 90.39039, 90.45312, 90.55574, 90.6293, 90.67559, 90.69638, 90.693535, 90.66931, 90.62608, 90.56623, 90.4921, 90.39684, 90.300255, 90.19653, 90.08777, 89.97542, 89.86078, 89.74513, 89.62964, 89.51496, 89.40164, 89.29024, 89.181206, 89.07475, 88.97101, 88.87012, 88.7721, 88.676605, 88.583206, 88.49145, 88.40098, 88.31178, 88.22392, 88.13745, 88.05242, 87.96885, 87.88672, 87.80605, 87.72684, 87.64909, 87.57282, 87.498055, 87.42471, 87.352455, 87.280876, 87.20955, 87.13802, 87.06573, 86.99203, 86.916306, 86.83819, 86.75831, 86.67755, 86.59681, 86.51706, 86.439674, 86.36613, 86.297905, 86.23633, 86.182144, 86.13594, 86.09829, 86.06955, 86.04905, 86.03585, 86.029015, 86.02752, 86.030045, 86.03515, 86.04142, 86.047516, 86.05247, 86.05541, 86.05548, 86.051994, 86.04503, 86.034904, 86.02192, 86.006424, 85.988914, 85.969955, 85.95009, 85.92979, 85.90921, 85.888405, 85.86741, 85.84625, 85.82488, 85.803215, 85.781166, 85.758644, 85.73551, 85.71162, 85.68681, 85.66099, 85.63419, 85.606544, 85.57815, 85.54914, 85.51978, 85.490364, 85.46119, 85.4325, 85.418365, 85.39047, 85.36306, 85.336105, 85.30956, 85.28338, 85.257515, 85.23192, 85.20665, 85.18189, 85.15551, 85.1325, 85.11056, 85.08974, 85.0701, 85.05169, 85.03451, 85.01852, 85.00367, 84.989914, 84.977234, 84.96566, 84.9552, 84.945885, 84.93753, 84.929794, 84.9223, 84.91468, 84.90646, 84.89706, 84.885864, 84.872314, 84.85601, 84.836784, 84.814476, 84.78892, 84.760025, 84.72775, 84.69209, 84.65301, 84.610435, 84.56428, 84.51442, 84.46076, 84.403305, 84.34214, 84.27738, 84.209145, 84.13766, 84.063324, 83.98653, 83.90767, 83.8273, 83.74617, 83.665, 83.58454, 83.5054, 83.428055, 83.35298, 83.28063, 83.21135, 83.14533, 83.082756, 83.02381, 82.96846, 82.91641, 82.867386, 82.82107, 82.77684, 82.73371, 82.690674, 82.646736, 82.6016, 82.55585, 82.51008, 82.46493, 82.42101, 82.37896, 82.33941, 82.30297, 82.26992, 82.240074, 82.22629, 82.200874, 82.17803, 82.15685, 82.13622, 82.11502, 82.09221, 82.06708, 82.03904, 82.007515, 81.97193, 81.93188, 81.88697, 81.83684, 81.78118, 81.72009, 81.653824, 81.58261, 81.50677, 81.427, 81.34419, 81.259186, 81.17281, 81.08575, 80.99861, 80.912, 80.82651, 80.74249, 80.66023, 80.580025, 80.50213, 80.426765, 80.35411, 80.28436, 80.21768, 80.15415, 80.093796, 80.036674, 79.982796, 79.9321, 79.88448, 79.83554, 79.79406, 79.75522, 79.7188, 79.68457, 79.65233, 79.621956, 79.59338, 79.56653, 79.54133, 79.5178, 79.49599, 79.47593, 79.45764, 79.44097, 79.42573, 79.41172, 79.39873, 79.38647, 79.37463, 79.36291, 79.35101, 79.338844, 79.326324, 79.3134, 79.30004, 79.28643, 79.27279, 79.25936, 79.24637, 79.233925, 79.22215, 79.211136, 79.20091, 79.19111, 79.18123, 79.17078, 79.15922, 79.14586, 79.12995, 79.11074, 79.08752, 79.05979, 79.027176, 78.98924, 78.94565, 78.89639, 78.84155, 78.78123, 78.71555, 78.64485, 78.5695, 78.489914, 78.40644, 78.31942, 78.229164, 78.13597, 78.04012, 77.94173, 77.84085, 77.73756, 77.63189, 77.52397, 77.413895, 77.30178, 77.18769, 77.07132, 76.95225, 76.83005, 76.70441, 76.57563, 76.44427, 76.31087, 76.176155, 76.042015, 75.91074, 75.78465, 75.66607, 75.55748, 75.461426, 75.380455, 75.31696, 75.2724, 75.24785, 75.24439, 75.262825, 75.30215, 75.36062, 75.436516, 75.52802, 75.63284, 75.74848, 75.87244, 76.00225, 76.135735, 76.27082, 76.40544, 76.5376, 76.665855, 76.78902, 76.905876, 77.0153, 77.12625, 77.218056, 77.30071, 77.37384, 77.43749, 77.49187, 77.537186, 77.573685, 77.60185, 77.622246, 77.63542, 77.64193, 77.64223, 77.636734, 77.62589, 77.61013, 77.58989, 77.565605, 77.537735, 77.50669, 77.47283, 77.43649, 77.39799, 77.35764, 77.31569, 77.27232, 77.22776, 77.18216, 77.135544, 77.087845, 77.03902, 76.98895, 76.93721, 76.883224, 76.82644, 76.766266, 76.701904, 76.63251, 76.55721, 76.47526, 76.386444, 76.2908, 76.18835, 76.079185, 75.96398, 75.8436, 75.7189, 75.590744, 75.45994, 75.327286, 75.19359, 75.059654, 74.92641, 74.79482, 74.66587, 74.540504, 74.419586, 74.303955, 74.19443, 74.09175, 73.9961, 73.90743, 73.82569, 73.75074, 73.68189, 73.618225, 73.55881, 73.502716, 73.44902, 73.39677, 73.34501, 73.29282, 73.239456, 73.21211, 73.15566, 73.0963, 73.03376, 72.968475, 72.90095, 72.83166, 72.761215, 72.69038, 72.61992, 72.585075, 72.51655, 72.44943, 72.38339, 72.318054, 72.25311, 72.188484, 72.12417, 72.060196, 71.99662, 71.927574, 71.86615, 71.806526, 71.749214, 71.69476, 71.64376, 71.59677, 71.5543, 71.51631, 71.48262, 71.45303, 71.4272, 71.40383, 71.38132, 71.358055, 71.332405, 71.302536, 71.26657, 71.222626, 71.16892, 71.13807, 71.067856, 70.98565, 70.89065, 70.7824, 70.66093, 70.52628, 70.37853, 70.2184, 70.04756, 69.867775, 69.77507, 69.58523, 69.39154, 69.19663, 69.00311, 68.81352, 68.62998, 68.454445, 68.28887, 68.13509, 67.99416, 67.92875, 67.808495, 67.70295, 67.61222, 67.53547, 67.471756, 67.42016, 67.37935, 67.347435, 67.32246, 67.302444, 67.28546, 67.26953, 67.25271, 67.23303, 67.20867, 67.17799, 67.13937, 67.09122, 67.03262, 66.96389, 66.8854, 66.797554, 66.701355, 66.59874, 66.49178, 66.382515, 66.27302, 66.16542, 66.06182, 65.96435, 65.874886, 65.79494, 65.725945, 65.66938, 65.62636, 65.59744, 65.58313, 65.58391, 65.59991, 65.63056, 65.67525, 65.70266, 65.76719, 65.84383, 65.931496, 66.0291, 66.135574, 66.25012, 66.372025, 66.50059, 66.63513, 66.7045, 66.84718, 66.99482, 67.14705, 67.303345, 67.46289, 67.62485, 67.78838, -999.0, -999.0, -999.0, -999.0, 68.530685, 68.69492, 68.85778, 69.01864, 69.17691, 69.33242, 69.48518, 69.63524, 69.70925, 69.855286, 69.94164, 70.083496, 70.2228, 70.359604, 70.49385, 70.625465, 70.75437, 70.88051, 71.00395, 71.124825, 71.24326, 71.3594, 71.4734, 71.585464, 71.695786, 71.804535, 71.91177, 72.01748, 72.121666, 72.22427, 72.324936, 72.42317, 72.51847, 72.61036, 72.69858, 72.78295, 72.86329, 72.939445, 73.011475, 73.07953, 73.14376, 73.174484, 73.23327, 73.28865, 73.340836, 73.39001, 73.436386, 73.48021, 73.521736, 73.5612, 73.59876, 73.63435, 73.66792, 73.69939, 73.72874, 73.75603, 73.78132, 73.80468, 73.82614, 73.84575, 73.863495, 73.87942, 73.89358, 73.90617, 73.91739, 73.92743, 73.936485, 73.944756, 73.95245, 73.95977, 73.96685, 73.97371, 73.98034, 73.986755, 73.99297, 73.99908, 74.00514, 74.01124, 74.01754, 74.02432, 74.031906, 74.0406, 74.04544, 74.05608, 74.067986, 74.08109, 74.095345, 74.110695, 74.12707, 74.14442, 74.16266, 74.18164, 74.201164, 74.22104, 74.24105, 74.26097, 74.280556, 74.29955, 74.31772, 74.334915, 74.35106, 74.36605, 74.381134, 74.39359, 74.40493, 74.415215, 74.424545, 74.43311, 74.44118, 74.448975, 74.45676, 74.46474, 74.47311, 74.48206, 74.49177, 74.50215, 74.51304, 74.52424, 74.53559, 74.54697, 74.55829, 74.56944, 74.580376, 74.591156, 74.596535, 74.607376, 74.61844, 74.62984, 74.6416, 74.65375, 74.66631, 74.67928, 74.69262, 74.70626, 74.720146, 74.73426, 74.74862, 74.76324, 74.77814, 74.793335, 74.80882, 74.82459, 74.840645, 74.85693, 74.87335, 74.88978, 74.90609, 74.92226, 74.93835, 74.95448, 74.97075, 74.98724, 75.00402, 75.02113, 75.038635, 75.056526, 75.07471, 75.09306, 75.11148, 75.129875, 75.14823, 75.16654, 75.18479, 75.202995, 75.221214, 75.23954, 75.248764, 75.26738, 75.286354, 75.30589, 75.32617, 75.34737, 75.369484, 75.392456, 75.41621, 75.440605, 75.4652, 75.48931, 75.51228, 75.53346, 75.55247, 75.56905, 75.58296, 75.594, 75.6024, 75.608635, 75.613174, 75.61648, 75.61872, 75.619896, 75.62003, 75.619125, 75.617226, 75.61441, 75.61073, 75.60626, 75.600945, 75.594635, 75.58723, 75.57858, 75.56859, 75.557144, 75.544136, 75.52945, 75.51292, 75.4923, 75.471115, 75.4474, 75.421326, 75.39321, 75.363396, 75.33222, 75.30013, 75.2676, 75.235115, 75.20321, 75.172745, 75.15838, 75.13202, 75.109695, 75.091934, 75.07834, 75.0684, 75.06161, 75.05767, 75.05667, 75.05875, 75.06402, 75.07261, 75.08461, 75.10011, 75.11921, 75.14165, 75.16657, 75.19304, 75.22009, 75.24698, 75.27327, 75.29859, 75.32255, 75.344826, 75.365234, 75.383575, 75.39968, 75.41338, 75.4246, 75.43323, 75.43918, 75.44245, 75.4432, 75.44163, 75.437904, 75.432236, 75.424835, 75.41593, 75.40574, 75.394455, 75.38225, 75.36927, 75.355675, 75.3416, 75.32717, 75.312485, 75.29766, 75.28279, 75.26793, 75.25312, 75.23842, 75.231125, 75.216606, 75.202156, 75.18773, 75.17326, 75.158676, 75.143845, 75.12866, 75.11301, 75.09681, 75.08002, 75.06258, 75.04446, 75.02578, 75.00678, 74.98772, 74.96879, 74.94989, 74.93073, 74.911, 74.89042, 74.87979, 74.85794, 74.8354, 74.81231, 74.78884, 74.76527, 74.741875, 74.71896, 74.69667, 74.674736, 74.65284, 74.630684, 74.607994, 74.58469, 74.56066, 74.53584, 74.51019, 74.483734, 74.45653, 74.42861, 74.40006, 74.37104, 74.341705, 74.31222, 74.28274, 74.253426, 74.22442, 74.19588, 74.167885, 74.14038, 74.11058, 74.08379, 74.05717, 74.030525, 74.00366, 73.976395, 73.94863, 73.92051, 73.8922, 73.86386, 73.83567, 73.8078, 73.78043, 73.753746, 73.72785, 73.70276, 73.67845, 73.65491, 73.6321, 73.60998, 73.58846, 73.56749, 73.5572, 73.53701, 73.51741, 73.49844, 73.48018, 73.46272, 73.44624, 73.43089, 73.416794, 73.40383, 73.3917, 73.3801, 73.36873, 73.3572, 73.34508, 73.33193, 73.31736, 73.301346, 73.28412, 73.26592, 73.246994, 73.22761, 73.20808, 73.18869, -999.0, -999.0, 73.13374, 73.11679, 73.10063, 73.0853, 73.07083, 73.057274, 73.05085, 73.03867, 73.02733, -999.0, -999.0, -999.0, -999.0, -999.0, 72.96976, 72.96526, 72.956184, 72.94691, 72.937325, 72.927345, 72.91697, 72.90629, 72.89537, 72.88429, 72.87306, 72.861664, 72.85589, 72.84417, 72.832275, 72.82038, 72.80873, 72.79754, 72.78696, 72.77691, 72.7673, 72.758026, 72.74897, 72.74446, 72.73538, 72.72606, 72.71631, 72.70598, 72.69497, 72.68316, 72.67044, 72.65677, -999.0, 72.62487, 72.60816, 72.59073, 72.572945, 72.5552, 72.53786, 72.52101, 72.50462, 72.488625, 72.47297, 72.457634, 72.45009, 72.43521, 72.42062, 72.40632, 72.39227, 72.37848, 72.364914, 72.3516, 72.3387, 72.32635, 72.31471, 72.30921, 72.298874, 72.2895, 72.28114, 72.27387, 72.26775, 72.262825, 72.25913, 72.256714, 72.25541, 72.25493, 72.254906, 72.25513, 72.255325, 72.25479, 72.252754, 72.248436, 72.24114, 72.23031, 72.2154, 72.19588, 72.184296, 72.158035, 72.12861, 72.09717, 72.06483, 72.03226, 71.999794, 71.96778, 71.936554, 71.90617, 71.87654, 71.847534, 71.81904, 71.790764, 71.76231, 71.73326, 71.70322, 71.67182, 71.63872, 71.60359, 71.56612, 71.546486, 71.50558, 71.46268, 71.41803, 71.37189, 71.32456, 71.276375, 71.22767, 71.1787, 71.12966, 71.08069, 71.03193, 70.983536, 70.93567, 70.8885, 70.84219, 70.79689, 70.7527, 70.70969, 70.667946, 70.62754, 70.58851, 70.550865, 70.51463, 70.47982, 70.446365, 70.41419, 70.38323, 70.35343, 70.324745, 70.29716, 70.28377, 70.257774, 70.23272, 70.208405, 70.18462, 70.1612, 70.138016, 70.115, 70.092094, 70.06925, 70.05782, 70.0349, 70.01178, 69.988365, 69.964615, 69.94074, 69.91701, 69.89367, 69.870926, 69.84878, 69.82505, 69.80401, 69.78341, 69.76315, 69.74312, 69.7232, 69.70331, 69.68342, 69.663506, 69.64356, 69.62354, 69.61348, 69.59319, 69.572624, 69.5517, 69.53044, 69.50898, 69.48744, 69.46594, 69.4445, 69.42313, 69.40179, 69.39112, 69.36978, 69.34833, 69.32666, 69.30467, 69.28227, 69.25942, 69.23609, 69.212234, 69.18788, 69.16313, 69.150665, 69.12561, 69.100525, 69.07551, 69.05059, 69.02583, 69.00128, 68.97704, 68.95324, 68.930016, 68.90751, 68.89654, 68.875206, 68.854675, 68.83498, 68.81611, 68.79811, 68.78099, 68.76477, 68.74945, 68.735, 68.72136, 68.714836, 68.70233, 68.69049, 68.67921, 68.66835, 68.65783, 68.64751, 68.63726, 68.62695, 68.61646, 68.60566, 68.59443, 68.582634, 68.57016, 68.557, 68.54321, 68.52886, 68.514046, 68.49905, 68.484375, 68.47053, 68.457985, 68.447044, 68.437836, 68.430466, 68.42503, 68.421326, 68.41882, 68.41701, 68.41537, 68.413536, 68.412476, 68.40993, 68.40662, 68.40233, 68.39691, 68.39023, 68.38214, 68.37258, 68.36179, 68.34885, 68.336426, 68.32365, 68.310616, 68.29743, 68.28419, 68.270966, 68.257805, 68.24471, 68.231735, 68.21888, 68.21252, 68.19992, 68.18754, 68.17539, 68.163445, 68.15162, 68.13983, 68.12799, 68.116035, 68.10391, 68.09156, 68.07893, 68.06589, 68.05225, 68.03784, 68.022484, 68.006256, 67.989395, 67.97216, 67.954796, 67.93753, 67.92899, 67.91224, 67.89608, 67.880615, 67.86573, 67.851234, 67.836945, 67.82287, 67.809525, 67.797585, 67.792336, 67.783676, 67.77761, 67.77406, 67.772964, 67.77419, 67.77707, 67.780426, 67.78309, 67.78389, 67.78187, 67.776276, 67.7719, -999.0, 67.741875, 67.71939, 67.6926, 67.66204, 67.62828, 67.5919, 67.55349, 67.51365, 67.47291, 67.43158, 67.38994, 67.34826, 67.306725, 67.26525, 67.22369, 67.18188, 67.13968, 67.09692, 67.07527, 67.03137, 66.98652, 66.9408, 66.89453, 66.84801, 66.801575, 66.75608, 66.71283, 66.67315, -999.0, 66.609184, 66.59677, 66.576385, 66.56209, 66.55377, 66.55032, 66.55038, 66.55255, 66.55575, 66.559845, 66.56498, 66.57128, 66.578865, 66.58772, -999.0, -999.0, -999.0, -999.0, 66.64905, 66.66345, 66.677956, 66.68658, 66.70059, 66.7139, 66.72617, 66.73694, 66.74558, 66.7515, 66.75411, 66.75314, 66.74862, 66.745026, 66.7352, 66.72204, 66.70627, 66.68873, 66.670265, 66.65161, 66.633156, 66.615204, 66.598076, 66.582, 66.566925, 66.55272, 66.539276, 66.52648, -999.0, -999.0, -999.0, -999.0, -999.0, 66.45737, 66.45167, 66.44003, 66.42817, -999.0, -999.0, -999.0, 66.38445, 66.3757, -999.0, -999.0, 66.35708, 66.353195, 66.35006, 66.347374, 66.34442, 66.34006, 66.333145, 66.32257, 66.30785, 66.289085, 66.26641, 66.23995, 66.20992, 66.1766, 66.14027, 66.10122, 66.05978, 66.016304, 65.97118, 65.92477, 65.87739, 65.82936, 65.78098, 65.75676, 65.708374, 65.660065, 65.61181, 65.563576}
u_wind =
  {0.7894132, -999.0, -999.0, 3.4071336, 3.9029899, -999.0, -999.0, -999.0, 4.6359396, 4.749648, 4.8832197, 5.0418286, 5.2131844, 5.3898425, 5.566017, 5.7351446, 5.893747, 6.038948, 6.168397, 6.2805977, 6.3749604, 6.452142, 6.5124655, 6.55603, 6.5830884, 6.5951996, 6.59435, 6.582454, 6.561498, 6.5331435, 6.4986887, 6.4598117, 6.4192495, 6.3799486, 6.343356, 6.309845, 6.2790384, 6.249219, 6.2190833, 6.1887193, 6.1583595, 6.128047, 6.097769, 6.0668244, 6.033945, 5.998526, 5.9610453, 5.921605, 5.879403, 5.8337193, 5.7861238, 5.739623, 5.6966023, 5.6586213, 5.6268897, 5.601078, 5.580619, 5.565464, 5.5556645, 5.551304, 5.553555, 5.563857, 5.586012, 5.62404, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 6.5163116, 6.5826406, 6.630386, 6.65151, -999.0, 6.6021576, -999.0, -999.0, -999.0, 6.1813374, -999.0, 5.8397374, -999.0, 5.4723816, -999.0, 5.1454525, 5.01422, 4.91174, -999.0, -999.0, -999.0, -999.0, -999.0, 4.85141, 4.9097095, 4.977366, 5.0479302, 5.1154385, 5.174975, 5.221947, 5.2533946, 5.2668567, 5.2615333, 5.237795, 5.196979, 5.1422043, 5.076575, 5.0036263, 4.927131, 4.8512063, 4.780157, 4.7181387, 4.6689897, 4.636502, 4.623251, 4.6317034, 4.66281, 4.717066, 4.7949686, 4.8963146, 5.0200453, 5.1625524, 5.3201528, 5.488454, 5.662737, 5.8381314, 6.009605, 6.172442, 6.322833, 6.4570475, 6.5727763, 6.6678405, 6.741679, 6.7945895, 6.828404, 6.847112, 6.8554177, 6.859749, 6.8662257, 6.8792925, 6.9032736, 6.9437823, 7.0068254, 7.096701, 7.215137, 7.3634377, 7.54107, 7.7472835, 7.9809694, 8.240527, 8.522248, 8.820094, 9.127767, 9.438577, 9.7462435, 10.047094, 10.366606, 10.643319, 10.903747, 11.144074, 11.359994, 11.548314, 11.709758, 11.845613, 11.958907, 12.053693, 12.134822, 12.208315, 12.280513, 12.35853, 12.449581, 12.560072, 12.696074, 12.861518, 13.058629, 13.289461, 13.55444, 13.853358, 14.18218, 14.535666, 14.905976, 15.284276, 15.665944, 16.049902, 16.431917, 16.801126, 17.146776, 17.463413, 17.746899, 17.99385, 18.203005, 18.373865, 18.508331, 18.608334, 18.675766, 18.712692, 18.721655, -999.0, 18.66723, 18.609838, 18.536, 18.446913, 18.343542, 18.22731, 18.099842, 17.963789, 17.823023, 17.681072, 17.540949, 17.405708, 17.278746, 17.16356, 17.063692, 16.982721, 16.923944, 16.889559, 16.881086, 16.897026, 16.93532, 16.993484, 17.068525, 17.156857, 17.254023, 17.355286, 17.45521, 17.548471, 17.630754, 17.697931, 17.745173, 17.767466, 17.761185, 17.725119, 17.657639, 17.556648, 17.42029, 17.250477, 17.051952, 16.832254, 16.601843, 16.367378, 16.125523, 15.872957, 15.615123, 15.360312, 15.114519, 14.882374, 14.667856, 14.473113, 14.300385, 14.152484, 14.032024, 13.93897, -999.0, 13.828338, 13.808262, 13.8097315, 13.829515, 13.863969, 13.908411, 13.957552, 14.010789, 14.052892, 14.084435, 14.1025, 14.104378, 14.088086, 14.051976, 13.995066, 13.916519, 13.81367, 13.682379, 13.521195, 13.336845, 13.137955, 12.9356165, 12.741115, 12.555214, 12.370098, 12.183723, 12.004246, 11.839903, 11.696023, 11.577193, 11.485972, 11.4236145, -999.0, 11.391067, -999.0, -999.0, 11.5789585, 11.695656, 11.834062, 11.986879, 12.14373, 12.297477, 12.447189, 12.591574, 12.724789, 12.839873, 12.931208, 12.994037, 13.024511, 13.020008, 12.978842, 12.90196, 12.790963, 12.648556, -999.0, 12.283833, 12.07185, 11.848381, 11.620787, 11.3965025, 11.182623, 10.986051, 10.812512, 10.666854, 10.553316, 10.475194, 10.435235, 10.434461, 10.473129, 10.548126, 10.654463, 10.786099, 10.935771, 11.095903, 11.258295, 11.414593, 11.55612, 11.674147, 11.76134, 11.811604, 11.819894, 11.783101, 11.698989, 11.568273, 11.392673, 11.175971, 10.9233055, 10.640782, 10.335838, 10.016453, 9.692021, 9.372176, 9.0661955, 8.783166, 8.531546, 8.319141, 8.152519, 8.035478, 7.9712973, 7.9625645, 8.011436, 8.117243, 8.232334, 8.427387, 8.667178, 8.946214, 9.258147, 9.596349, 9.955181, 10.368033, 10.754787, 11.147484, 11.540675, 11.926601, 12.297276, 12.646156, 12.96718, 13.254226, 13.501785, 13.704648, 13.859632, 13.963473, 14.013899, 14.009048, 13.948647, 13.83483, 13.670304, 13.461564, 13.215045, 12.9391775, 12.643255, 12.338267, 12.036704, 11.7507, 11.491182, 11.268893, 11.090961, 10.964678, 10.895691, 10.888068, 10.941948, 11.051519, 11.21095, 11.411497, 11.644176, 11.898734, 12.164131, 12.427839, 12.676266, 12.8971405, 13.081189, 13.219359, 13.306412, 13.338109, 13.314224, 13.237031, 13.109566, 12.936978, 12.725071, 12.481963, 12.216079, 11.936106, 11.650911, 11.368674, 11.096767, 10.841804, 10.608292, 10.400546, 10.221134, 10.071947, 9.953032, 9.8633175, 9.8026085, 9.7712555, 9.768959, 9.793555, 9.842796, 9.914934, 10.008059, 10.1191, 10.24481, 10.385202, 10.544577, 10.724991, 10.916605, 11.107245, 11.293131, 11.47527, 11.652718, 11.8233, 11.984784, 12.1340065, 12.267648, 12.38425, 12.483261, 12.563642, 12.624893, 12.667028, 12.69198, -999.0, 12.697636, 12.6783285, 12.648776, 12.609363, 12.562027, 12.509342, 12.453603, 12.396135, 12.338192, 12.281954, 12.229907, 12.184006, 12.146452, 12.120273, 12.110131, 12.12072, 12.153899, 12.210738, 12.293022, 12.402282, 12.539666, 12.704611, 12.896748, 13.114248, 13.355049, -999.0, 13.893574, 14.182236, 14.475628, 14.767603, 15.051101, 15.318877, 15.563069, 15.775001, 15.945237, 16.065046, 16.126879, 16.131084, 16.078703, 15.973854, 15.821369, 15.622691, 15.378105, 15.091702, 14.775707, 14.441802, 14.100966, 13.764822, 13.443438, 13.145678, 12.879901, 12.6513605, 12.4654455, -999.0, 12.221082, 12.158985, 12.131703, 12.133758, 12.157166, 12.194344, 12.2378845, 12.279756, 12.312324, 12.3279, 12.321435, 12.290341, 12.232437, 12.148933, 12.040963, 11.912222, 11.766703, 11.609397, 11.446234, 11.283725, 11.129108, 10.989552, 10.869891, 10.7752, 10.707883, 10.669467, 10.66063, 10.680183, 10.726694, 10.796316, 10.885128, 10.987897, 11.098965, 11.21285, 11.324061, 11.427283, 11.517776, 11.590274, 11.640472, 11.664037, 11.660055, 11.629049, 11.571737, 11.490473, 11.388127, 11.269539, 11.139041, 11.000761, 10.859334, 10.72225, 10.598668, 10.495535, 10.415696, 10.362624, 10.337748, 10.3420725, 10.374447, 10.432317, 10.512739, 10.622309, 10.736759, -999.0, 10.991447, 11.1228075, 11.250696, 11.372705, 11.48802, 11.595811, 11.696686, 11.791664, 11.883392, 11.974874, 12.068281, 12.165596, 12.26774, 12.374095, 12.483766, 12.594348, 12.703281, 12.806781, 12.900592, 12.979907, 13.039418, 13.074217, 13.080429, 13.054558, 12.995928, 12.904352, 12.782216, 12.633591, 12.465008, 12.286201, 12.106897, 11.937429, 11.7883005, 11.669731, 11.591831, 11.563202, 11.590904, 11.679942, 11.830963, 12.043796, 12.314478, 12.6379595, 13.006898, 13.412622, 13.84696, 14.301938, 14.76918, 15.239621, 15.704261, 16.155947, 16.5884, 16.997463, 17.381166, 17.737413, 18.064457, 18.360697, 18.62518, 18.857094, 19.055485, 19.219322, 19.347702, 19.439787, 19.494732, 19.511238, 19.48781, 19.422245, 19.311989, 19.155317, 18.951685, 18.70091, 18.404703, 18.064987, 17.684643, 17.266977, 16.815918, 16.336348, 15.833965, 15.316249, 14.790523, 14.263381, 13.741542, 13.232707, 12.745016, 12.285706, 11.860606, 11.475096, 11.132706, 10.836866, 10.591563, 10.384799, 10.256347, 10.184575, 10.1681385, 10.203185, 10.286519, 10.416485, 10.591255, 10.805681, 11.053096, 11.327398, 11.622555, 11.932432, 12.250938, 12.571997, 12.890298, 13.2008505, 13.499452, 13.782887, 14.048589, 14.296103, 14.525282, 14.737687, 14.935347, 15.120696, 15.296776, 15.467251, 15.6367235, 15.809689, 15.989474, 16.179192, 16.380196, 16.59291, 16.817608, 17.0538, 17.300592, 17.555866, 17.81746, 18.083422, 18.351717, 18.619953, 18.885654, 19.146969, 19.402903, 19.652184, 19.892275, 20.120493, 20.334345, 20.531378, 20.709251, 20.865099, 20.995571, 21.094912, 21.155972, 21.171165, 21.133932, 21.046974, 20.920965, 20.760725, 20.560843, 20.315895, 20.026398, 19.694138, 19.327156, 18.939245, 18.542164, 18.146374, 17.76294, 17.40174, 17.072655, 16.783195, 16.539154, 16.344255, 16.197676, 16.098661, 16.042404, 16.023573, 16.033253, 16.060858, 16.0953, 16.124544, 16.136923, 16.122778, 16.07235, 15.979335, 15.838081, 15.645721, 15.402073, 15.108728, 14.772416, 14.400357, 14.004361, 13.59719, 13.192951, 12.806646, 12.452029, 12.141088, 11.884842, 11.689978, 11.563333, 11.508201, 11.526366, 11.625473, 11.776397, 11.971256, 12.19329, 12.431636, 12.687178, 12.958777, 13.230053, 13.480975, 13.700194, 13.88252, 14.0257225, 14.133973, 14.210432, 14.254109, 14.263789, 14.242517, -999.0, 14.130736, 14.057686, 13.984452, 13.913815, 13.847907, 13.788105, 13.7351675, 13.688577, -999.0, 13.608912, 13.574664, 13.543961, 13.516695, 13.492633, 13.470503, 13.448552, 13.42632, 13.404878, 13.385162, 13.367809, 13.353609, 13.344237, 13.341593, 13.346131, 13.3569975, 13.373411, 13.394526, 13.41941, 13.446328, 13.473051, 13.495007, 13.505975, 13.500556, -999.0, 13.4527855, 13.389947, 13.300574, 13.184656, 13.04497, 12.884222, 12.704433, 12.5078335, 12.299891, 12.08841, 11.882408, 11.692295, 11.526379, 11.385673, 11.27022, 11.182406, 11.125315, 11.101252, 11.111666, 11.1570215, 11.2351465, 11.343898, 11.481548, 11.645758, 11.829187, 12.020905, 12.214113, 12.408257, 12.601052, 12.7842865, -999.0, 13.097034, 13.230904, 13.352525, 13.460988, 13.557203, 13.64769, 13.739314, 13.835724, 13.939785, 14.056574, 14.192229, 14.350998, 14.53111, 14.729924, 14.943288, 15.166644, 15.39918, 15.6422825, 15.893095, 16.167929, 16.411358, 16.652029, 16.89277, 17.124851, 17.335217, 17.517159, 17.66988, 17.79158, -999.0, 17.948215, 17.991524, 18.020071, 18.038168, 18.049215, 18.058495, 18.073656, 18.101847, 18.147009, -999.0, 18.302044, 18.417852, 18.56135, 18.730972, 18.92415, 19.13461, 19.356098, 19.584486, 19.815866, 20.04342, 20.258238, 20.45299, 20.623388, -999.0, 20.87399, 20.946579, 20.98149, 20.979038, 20.94003, 20.86721, 20.763784, 20.634975, 20.486357, 20.323988, 20.154411, 19.984604, 19.821823, 19.672583, 19.541296, 19.432375, 19.349876, 19.297638, 19.27807, 19.291912, 19.338324, 19.412977, 19.511631, 19.630339, 19.764849, 19.910143, 20.061222, 20.215307, 20.371666, 20.527525, 20.675724, 20.80941, 20.927034, 21.028675, -999.0, 21.181252, -999.0, 21.266918, 21.28807, 21.296976, 21.29516, 21.282991, 21.260418, 21.2294, 21.194147, -999.0, 21.119844, 21.08055, 21.042274, 21.008366, 20.981045, 20.961563, 20.950926, -999.0, 20.957447, 20.976074, 21.00661, 21.04956, 21.104486, -999.0, 21.241463, 21.315258, 21.387554, 21.454874, 21.515099, 21.566927, 21.608677, 21.638536, 21.655655, 21.65561, 21.63925, 21.605774, 21.554916, 21.489147, 21.412958, 21.329498, 21.240044, 21.145649, 21.047205, 20.94591, 20.845726, 20.751848, 20.667265, 20.592464, 20.52789, 20.473595, 20.429964, 20.399206, 20.38397, 20.38436, 20.398233, -999.0, 20.45793, 20.498451, 20.542952, 20.589699, 20.63949, 20.694622, 20.755302, -999.0, 20.883831, 20.948679, 21.01219, 21.07113, 21.121506, 21.160355, 21.186062, -999.0, -999.0, 21.192604, 21.175018, 21.145184, 21.10185, 21.044413, 20.972906, 20.892174, 20.808802, 20.72629, 20.646524, 20.574053, 20.516766, 20.481398, 20.467018, 20.47111, 20.493776, 20.535704, 20.595757, -999.0, 20.755909, 20.85019, 20.950457, -999.0, -999.0, 21.242125, 21.31861, 21.376284, 21.413458, 21.428743, 21.421001, 21.389248, 21.331991, 21.247578, 21.135084, 20.99647, 20.83467, 20.656866, 20.471046, 20.282236, 20.094093, 19.91115, 19.738344, 19.580326, 19.440878, 19.323954, 19.233044, 19.17107, -999.0, 19.133108, 19.152632, 19.194551, 19.255934, 19.331654, 19.415886, 19.503466, 19.58963, 19.669939, 19.740765, 19.798243, 19.838476, 19.857805, 19.85459, 19.828152, 19.777168, 19.700401, 19.596956, 19.468922, 19.319187, 19.15447, 18.983131, 18.811686, 18.644716, 18.469631, 18.31765, 18.173254, 18.041567, 17.928125, 17.834412, 17.760134, -999.0, 17.664331, 17.636734, 17.617756, 17.603373, 17.588829, 17.569208, 17.54074, 17.499783, 17.43974, 17.35244, 17.231033, 17.081251, -999.0, 16.823795, 16.644966, -999.0, 16.294044, 16.10834, 15.919041, 15.741941, 15.587432, 15.4593935, 15.36252, 15.299965, 15.274238, 15.2876835, 15.342174, 15.438253, 15.574643, 15.752318, -999.0, 16.228378, 16.512314, 16.80641, 17.096067, 17.36723, 17.6089, 17.818434, 17.992035, 18.121527, 18.1983, 18.219198, 18.18474, 18.095821, 17.957731, 17.776575, 17.563814, 17.332111, -999.0, 16.865232, 16.65586, 16.476444, 16.336405, 16.241587, 16.197634, 16.208445, 16.277355, 16.405472, 16.590534, 16.826916, 17.101284, 17.400549, -999.0, 18.028044, 18.33409, 18.621044, 18.878574, 19.097078, 19.266602, 19.379927, 19.43101, 19.422344, 19.359673, 19.246838, 19.08796, 18.888653, 18.658964, 18.409954, 18.155481, 17.910267, 17.68436, 17.483982, 17.313286, 17.171436, 17.058422, 16.975773, 16.925203, 16.905413, 16.913183, 16.942205, -999.0, 17.024757, 17.06445, 17.095753, -999.0, 17.115692, 17.102808, 17.068449, 17.01145, 16.932491, 16.833055, 16.715565, 16.58402, 16.443434, 16.30057, 16.161737, 16.030102, 15.908444, 15.8001375, 15.708427, 15.636, 15.584188, 15.553913, 15.543836, 15.552435, 15.57832, 15.619903, 15.674946, 15.740495, 15.813604, 15.891076, -999.0, 16.0468, 16.11892, 16.182161, 16.232561, 16.268522, 16.291956, 16.303724, 16.302422, 16.286648, 16.257912, 16.219141, 16.1739, 16.126432, 16.079264, 16.031721, 15.983808, 15.9401455, 15.906472, -999.0, 15.8786545, 15.88572, 15.90551, 15.936375, 15.975268, 16.018885, 16.065283, 16.11308, 16.159824, -999.0, 16.23695, 16.261953, 16.275465, 16.278412, 16.272455, 16.256372, 16.227396, 16.185747, 16.136826, 16.085415, 16.031696, 15.974859, 15.914505, 15.85025, 15.783073, 15.716075, 15.651855, 15.591261, 15.53491, 15.483534, 15.4379015, 15.39957, 15.370677, 15.352431, 15.3438225, -999.0, 15.347425, 15.361273, 15.383934, 15.413243, 15.447319, 15.486837, 15.533154, 15.58496, 15.638465, 15.690293, 15.743057, 15.785953, 15.82628, 15.866674, 15.906525, 15.9439335, 15.979086, 16.01369, 16.048267, 16.080421, -999.0, 16.128983, 16.144089, 16.153143, 16.157043, 16.155813, 16.148182, 16.13341, 16.11262, 16.087008, 16.055302, 16.014977, 15.965491, 15.908756, 15.845885, 15.775833, -999.0, 15.610844, 15.5168705, 15.4169, 15.312551, 15.203533, 15.086563, 14.959528, 14.827654, 14.697656, 14.569648, 14.439981, 14.309545, 14.185629, 14.074028, 13.974879, 13.887786, 13.81556, 13.762283, -999.0, 13.723564, 13.742541, 13.788859, 13.862346, -999.0, 14.007075, 14.113899, 14.226099, 14.34258, 14.45836, 14.567028, 14.66343, 14.743742, 14.804152, 14.843124, 14.859223, -999.0, 14.824265, 14.777056, 14.714961, 14.64144, 14.559226, 14.47126, 14.380414, 14.289247, 14.199528, 14.112944, 14.032818, 13.963404, -999.0, 13.86633, 13.834498, 13.808615, 13.783275, 13.755399, 13.724287, 13.688388, 13.645316, 13.592434, -999.0, 13.449162, 13.356455, 13.250997, 13.134459, 13.011788, 12.888231, -999.0, 12.712727, 12.609882, 12.52274, 12.455459, 12.411304, 12.392805, 12.39921, 12.426415, 12.471659, 12.53274, 12.615233, 12.699389, 12.78729, -999.0, 12.951925, -999.0, 13.06568, 13.092568, 13.096258, 13.074479, 13.026005, 12.950661, 12.850728, 12.729596, 12.587116, 12.419395, 12.224057, 12.00737, 11.77691, 11.538162, 11.296512, 11.057022, 10.821679, 10.590637, 10.36078, 10.128857, 9.899735, 9.682283, 9.485431, -999.0, 9.174188, 9.0484705, -999.0, 8.820043, 8.725564, 8.646145, 8.580267, 8.526752, 8.482984, 8.445874, 8.411641, 8.376226, 8.33842, 8.298532, 8.257043, -999.0, 8.174874, 8.1358185, 8.098813, 8.064625, 8.033997, 8.007607, -999.0, 7.9702373, 7.960613, -999.0, 7.962552, 7.975053, 7.9957995, 8.025021, 8.062584, 8.107248, 8.157369, 8.21055, 8.264344, 8.318405, 8.373281, 8.429578, -999.0, 8.548365, 8.608913, 8.6682, 8.727177, 8.787437, 8.850501, 8.917788, 8.9891205, 9.062176, 9.136031, 9.211963, -999.0, 9.369848, 9.443517, 9.50793, 9.559654, 9.59579, 9.615547, 9.617942, 9.60202, 9.567029, 9.513895, -999.0, 9.405904, 9.319842, 9.227559, 9.133658, 9.042704, 8.958174, 8.88068, 8.810952, 8.750002, 8.698617, 8.652734, 8.6196575, 8.594389, 8.576841, 8.566512, 8.561868, 8.561323, 8.563735, -999.0, 8.573507, 8.57951, 8.585563, 8.591633, 8.597681, 8.604531, -999.0, 8.626671, 8.647244, 8.676871, 8.715642, 8.763864, 8.821954, 8.890349, 8.969177, -999.0, 9.157211, 9.264427, 9.378441, 9.497328, 9.619262, 9.743593, 9.870143, 9.998969, 10.130024, 10.261449, 10.388992, 10.509407, 10.623343, 10.7318325, 10.8346615, 10.9314375, 11.022348, 11.108065, 11.189346, 11.266636, 11.339973, 11.407516, 11.466939, 11.517814, 11.561073, 11.597145, 11.626062, 11.647954, 11.663414, 11.673131, 11.67816, 11.679837, 11.679551, 11.678972, 11.679859, -999.0, 11.695068, 11.714256, 11.744531, 11.787519, 11.843456, 11.911671, 11.989316, 12.074064, 12.165737, 12.264322, -999.0, 12.417104, 12.51413, 12.6028, 12.680237, 12.74548, 12.800369, 12.846376, 12.885661, 12.9205065, 12.954296, 12.990754, 13.0339985, 13.088777, 13.159905, 13.252112, 13.371364, 13.521632, 13.705603, 13.918089, 14.149876, 14.397986, 14.664872, 14.950447, 15.247023, 15.546481, 15.8410635, 16.122269, 16.382864, 16.617878, 16.82265, 16.995214, 17.13282, 17.233477, -999.0, 17.323427, 17.32179, 17.295643, 17.247997, 17.182144, 17.100584, 17.005213, 16.885422, 16.763988, 16.635145, 16.505714, 16.379766, 16.258606, 16.144707, 16.045774, 15.970429, 15.925848, 15.91876, 15.95456, 16.03504, 16.160297, 16.325335, 16.525724, 16.76195, 17.035086, 17.338884, 17.66202, 17.998396, 18.348701, 18.71152, 19.075031, 19.425554, 19.754515, 20.055805, 20.32348, -999.0, 20.743761, 20.890198, 20.990505, 21.042706, 21.045319, 20.998167, -999.0, 20.766111, 20.59112, 20.385256, 20.155056, 19.907589, 19.651594, 19.397236, 19.154047, 18.930056, 18.733349, 18.569958, 18.44554, 18.364107, 18.328135, 18.339077, 18.395094, 18.493967, 18.629671, 18.795547, 18.98376, 19.185686, 19.39324, 19.59886, 19.794798, 19.974434, 20.131023, 20.260782, 20.3609, 20.431152, 20.474106, 20.492342, 20.489697, 20.470133, 20.43727, 20.395016, 20.34658, 20.294317, 20.23851, 20.176153, 20.104937, 20.02286, 19.927698, 19.816221, 19.68466, 19.529322, 19.34718, 19.136364, 18.899734, 18.639801, 18.360922, 18.068203, 17.768675, 17.471079, 17.183817, 16.915041, 16.673391, 16.465694, 16.298956, 16.177515, 16.103819, 16.078373, 16.098463, 16.16237, 16.269428, 16.420366, 16.613895, 16.871655, 17.132544, 17.399288, 17.663017, 17.927378, 18.193075, 18.45436, 18.705458, 18.939596, 19.148827, 19.326618, 19.468075, 19.568193, 19.6245, 19.634764, 19.600466, -999.0, 19.410961, 19.265324, 19.091085, 18.89119, 18.670794, 18.442589, 18.219954, 18.012669, 17.829325, 17.677958, 17.565374, 17.498308, 17.482359, 17.522661, 17.620531, 17.775816, -999.0, 18.240582, 18.536362, 18.86467, 19.218912, 19.593939, 19.984455, 20.38041, 20.768913, 21.134329, 21.458878, 21.729788, 21.947424, 22.11342, -999.0, 22.301495, -999.0, 22.320772, 22.273565, 22.189222, 22.070158, 21.929749, 21.784113, 21.647837, -999.0, 21.452806, 21.404816, 21.392515, -999.0, 21.475838, 21.57161, 21.70327, 21.866896, -999.0, 22.257353, 22.46651, 22.67327, 22.873198, -999.0, -999.0, 23.30719, 23.42987, 23.518438, 23.576324, 23.60709, 23.615677, 23.605524, 23.57679, 23.52985, -999.0, 23.43207, 23.35434, -999.0, 23.18991, 23.109324, 23.03142, 22.959377, -999.0, 22.847994, 22.811241, 22.786125, 22.779943, -999.0, 22.822512, 22.870886, 22.939999, 23.035337, 23.160234, 23.31278, 23.49044, 23.689339, -999.0, 24.135136, 24.377533, 24.627249, 24.87569, 25.118347, 25.361717, 25.61101, -999.0, 25.956842, 26.135239, 26.264166, -999.0, 26.380903, 26.384983, 26.360973, 26.307852, 26.225702, 26.1184, -999.0, 25.923899, 25.789457, -999.0, 25.556664, 25.468227, -999.0, 25.35887, 25.340282, 25.347599, 25.380507, -999.0, 25.467741, 25.54105, 25.614073, -999.0, -999.0, 25.762365, 25.776855, 25.766241, 25.725374, 25.649115, 25.534935, 25.386158, 25.206621, -999.0, 24.767303, 24.518158, -999.0, -999.0, 23.777561, -999.0, 23.397879, 23.265991, 23.180809, 23.147503, 23.166489, 23.231236, 23.333496, 23.461557, -999.0, 23.759073, 23.926846, -999.0, 24.286129, 24.464117, 24.630114, 24.775164, 24.890833, 24.969387, 25.010553, -999.0, -999.0, -999.0, 24.954376, 24.910355, 24.865717, 24.826021, 24.795774, 24.779556, 24.782013, 24.807503, 24.85728, -999.0, -999.0, 25.074682, 25.18749, 25.311033, 25.446426, 25.59087, 25.734488, 25.86803, -999.0, -999.0, -999.0, 26.244368, 26.33512, -999.0, 26.515759, -999.0, 26.729963, 26.863522, 27.011497, -999.0, 27.246796, -999.0, 27.481941, 27.605906, 27.705349, 27.7739, 27.804886, -999.0, 27.737152, -999.0, 27.496866, 27.322779, -999.0, 26.87438, 26.601217, -999.0, 25.991901, 25.665792, 25.328108, 24.98182, 24.631418, 24.291794, 23.988474, 23.736511, 23.522606, 23.331068, 23.15643, 22.996557, 22.852491, 22.728561, 22.626308, 22.54249, -999.0, 22.447596, 22.409218, 22.393587, -999.0, 22.426945, 22.4766, 22.55091, -999.0, 22.778667, 22.931307, 23.103697, -999.0, 23.487354, 23.689888, 23.888817, 24.072754, 24.235895, 24.37888, 24.500898, 24.596848, 24.661549, 24.693554, 24.693283, 24.667439, -999.0, 24.588585, 24.56058, 24.559034, -999.0, 24.67589, 24.807732, 24.98821, 25.214264, -999.0, -999.0, 26.109503, 26.45742, 26.822628, 27.203667, 27.585232, -999.0, 28.096952, 28.364096, 28.55238, 28.657455, -999.0, -999.0, 28.575876, 28.450556, -999.0, 28.114288, 27.921917, 27.722376, 27.52323, 27.334703, 27.166195, 27.021908, 26.904259, 26.812023, 26.7416, 26.689528, 26.649633, 26.626663, -999.0, 26.618795, 26.632912, 26.657171, 26.69134, 26.736242, 26.793959, 26.868732, 26.963816, 27.07754, 27.207193, -999.0, 27.513922, 27.6887, 27.868338, 28.046785, 28.225698, 28.406548, 28.579672, -999.0, 28.795813, 28.904097, 28.98444, 29.040565, 29.077785, 29.099945, 29.109102, 29.107754, 29.09985, 29.089455, 29.07973, 29.073416, 29.071955, -999.0, 29.084064, 29.095577, -999.0, 29.12089, 29.13135, 29.136953, 29.134155, 29.11993, 29.09202, 29.0486, 28.989063, 28.913446, 28.824942, 28.728264, 28.628319, 28.530188, 28.435926, -999.0, 28.238892, 28.131088, -999.0, 27.904013, 27.787767, 27.672905, 27.5643, 27.466465, -999.0, -999.0, -999.0, -999.0, -999.0, 27.168861, -999.0, 27.147598, 27.15215, -999.0, 27.187366, 27.213968, 27.243979, 27.275663, -999.0, -999.0, 27.375624, 27.405638, -999.0, -999.0, 27.463934, 27.472448, 27.47303, 27.465462, -999.0, 27.431065, 27.407646, -999.0, 27.358591, 27.337358, 27.31903, 27.302235, 27.28534, 27.266378, 27.244009, -999.0, 27.191843, 27.161846, 27.127068, 27.086445, 27.0397, 26.979965, -999.0, 26.838778, -999.0, 26.668488, 26.586689, -999.0, 26.463524, 26.429861, 26.417692, 26.428205, -999.0, 26.487076, -999.0, 26.632587, 26.730375, -999.0, 26.970427, 27.100824, 27.229742, 27.352491, 27.441317, 27.54933, -999.0, 27.74803, 27.829556, 27.894903, 27.945097, 27.981207, 28.004961, 28.018215, 28.022505, 28.019308, -999.0, 27.996744, 27.980553, 27.962969, 27.94482, 27.925266, 27.903307, 27.880833, 27.86147, -999.0, 27.84056, 27.842302, 27.855995, 27.884613, 27.92792, -999.0, 28.050758, 28.125683, -999.0, 28.303114, 28.412928, 28.5336, -999.0, 28.779802, 28.890625, 28.985071, -999.0, 29.125158, -999.0, -999.0, -999.0, -999.0, -999.0, 29.189468, 29.163229, 29.131863, 29.09946, -999.0, 29.045204, 29.0291, -999.0, 29.031467, 29.052341, 29.085701, -999.0, 29.188908, 29.257908, -999.0, 29.421032, 29.507082, -999.0, 29.625885, 29.694166, 29.75254, 29.802223, -999.0, 29.884304, 29.917557, 29.94564, -999.0, 29.989948, 30.009144, 30.02924, 30.052023, -999.0, -999.0, 30.148579, -999.0, 30.244244, 30.30416, 30.36888, 30.432577, 30.492027, 30.54682, 30.596079, 30.638468, 30.67275, 30.698576, 30.71611, -999.0, 30.73198, 30.734015, -999.0, 30.72658, 30.715956, 30.698818, 30.67356, 30.638552, -999.0, 30.537931, 30.47478, 30.406895, 30.336824, 30.26274, 30.18173, 30.09549, 30.00937, -999.0, -999.0, 29.797281, 29.76092, 29.753742, -999.0, 29.798676, -999.0, -999.0, -999.0, 30.19129, -999.0, -999.0, 30.656996, 30.804895, 30.937843, -999.0, -999.0, -999.0, 31.315138, 31.375578, 31.419256, 31.446075, 31.456879, 31.456047, 31.448946, 31.435595, 31.411222, -999.0, -999.0, 31.24593, 31.157705, -999.0, 30.933891, 30.799814, 30.652323, -999.0, -999.0, 30.246443, 30.08498, -999.0, -999.0, 29.699303, -999.0, 29.583702, 29.577223, -999.0, 29.625387, 29.697178, 29.804192, 29.946835, -999.0, 30.322416, 30.533272, -999.0, 30.95704, -999.0, -999.0, 31.497528, 31.677782, 31.819542, 31.915268, -999.0, 31.947447, 31.87699, 31.747513, -999.0, -999.0, -999.0, 30.923939, 30.639385, 30.356722, 30.079466, 29.809507, -999.0, 29.336424, -999.0, 29.029785, 28.9459, 28.915316, -999.0, -999.0, 29.0423, 29.152397, 29.279371, 29.410263, 29.534685, 29.644054, 29.741539, -999.0, -999.0, -999.0, 30.010862, -999.0, 30.050915, 30.029984, -999.0, 29.92273, 29.84311, -999.0, -999.0, 29.588413, -999.0, 29.334661, 29.199017, -999.0, 28.942951, 28.832075, -999.0, 28.638512, -999.0, -999.0, 28.453651, 28.410461, 28.393616, 28.40243, 28.43628, 28.493603, -999.0, -999.0, -999.0, -999.0, 28.939089, 29.055573, 29.171865, 29.284103, 29.387388, 29.47674, -999.0, 29.60267, 29.644852, 29.67583, 29.695704, 29.70456, 29.702433, 29.689417, -999.0, 29.641537, 29.61311, 29.586527, -999.0, 29.553703, -999.0, 29.56258, 29.591812, 29.642601, 29.71349, 29.803053, 29.910841, 30.037022, 30.183294, 30.351639, 30.539587, 30.738678, -999.0, 31.149586, -999.0, -999.0, 31.715673, -999.0, 31.953077, 32.014717, 32.03727, 32.020172, 31.961641, 31.860376, 31.719038, -999.0, 31.330866, 31.084566, 30.802448, 30.492239, -999.0, -999.0, 29.711681, 29.477148, 29.300848, 29.177822, 29.109093, 29.094984, 29.132904, 29.218279, 29.349138, -999.0, 29.628876, 29.86021, 30.102266, 30.333914, -999.0, -999.0, -999.0, 31.055422, 31.186504, 31.294483, 31.383581, -999.0, 31.478819, 31.506737, 31.53246, 31.558666, 31.585758, 31.619032, 31.668089, 31.73905, -999.0, 31.875494, 31.97757, 32.082287, 32.18623, 32.291843, 32.401546, 32.510193, -999.0, -999.0, -999.0, -999.0, 32.87093, -999.0, 32.976566, 33.02664, 33.08101, -999.0, 33.20535, 33.276432, 33.35485, -999.0, -999.0, 33.601364, 33.733536, 33.894905, 34.08827, 34.308243, 34.5473, 34.794834, 35.041916, 35.29502, 35.567028, -999.0, -999.0, -999.0, 36.57007, 36.815666, 37.023796, 37.191307, 37.313942, -999.0, -999.0, -999.0, -999.0, 37.331806, 37.24202, -999.0, 36.996727, 36.853752, 36.706097, 36.55994, -999.0, 36.30223, 36.206593, -999.0, 36.088966, 36.064896, 36.065228, 36.089382, 36.133305, 36.192963, 36.26638, 36.352238, 36.44991, 36.55902, -999.0, 36.796482, 36.912907, 37.025326, 37.133682, 37.23714, 37.335114, -999.0, -999.0, -999.0, 37.6336, 37.700138, 37.755466, 37.802036, 37.841614, 37.874153, -999.0, 37.918865, 37.933247, 37.944714, 37.951912, 37.955963, -999.0, 37.948547, 37.935356, 37.915737, -999.0, 37.865364, 37.841408, -999.0, 37.8186, -999.0, 37.83757, 37.874683, 37.925644, 37.987793, -999.0, 38.159496, -999.0, 38.39183, -999.0, 38.638832, 38.748863, -999.0, -999.0, -999.0, 39.053513, 39.09525, 39.126526, 39.148827, -999.0, 39.16717, 39.17224, 39.17625, -999.0, 39.197, -999.0, 39.259182, 39.313217, -999.0, -999.0, 39.490005, 39.5644, 39.640133, 39.719578, -999.0, -999.0, 39.99943, -999.0, -999.0, 40.247967, -999.0, -999.0, 40.368114, 40.392, -999.0, -999.0, 40.407375, 40.401608, 40.393887, 40.38612, 40.38109, 40.382065, -999.0, 40.422096, 40.47065, -999.0, -999.0, -999.0, 40.848114, -999.0, 41.10853, -999.0, 41.3303, 41.489998, -999.0, 41.797176, -999.0, 42.016502, 42.08032, 42.1133, -999.0, 42.09358, -999.0, -999.0, -999.0, 41.81649, 41.689396, 41.551666, 41.412308, -999.0, -999.0, -999.0, 40.983936, 40.916798, -999.0, 40.839584, -999.0, 40.842583, 40.873707, 40.923756, -999.0, 41.066837, 41.150993, -999.0, 41.287937, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 41.69665, 41.70962, -999.0, 41.702805, -999.0, -999.0, 41.621433, 41.581654, 41.54163, -999.0, 41.48347, -999.0, 41.461273, 41.463867, -999.0, -999.0, 41.518337, -999.0, 41.57316, 41.60686, -999.0, 41.682137, 41.71801, -999.0, 41.757507, 41.770554, -999.0, 41.755177, 41.72184, -999.0, -999.0, -999.0, 41.430267, -999.0, 41.217, 41.095726, 40.97726, 40.898445, 40.901222, -999.0, -999.0, -999.0, 41.693863, -999.0, 41.795094, -999.0, 38.580704, -999.0, -999.0, -999.0, -999.0, -999.0, 4.675371, 1.1835966, -0.7451929, -999.0, -999.0, -999.0, -999.0, -0.9107407, -0.22643878, -999.0}
v_wind =
  {2.5820198, -999.0, -999.0, 12.137266, 13.843243, -999.0, -999.0, -999.0, 15.718887, 15.84257, 16.020079, 16.269403, 16.541306, 16.809044, 17.058474, 17.27197, 17.443542, 17.57014, 17.651833, 17.692045, 17.694344, 17.663286, 17.603897, 17.522234, 17.424559, 17.317402, 17.20749, 17.100801, 17.002377, 16.916975, 16.847118, 16.795055, 16.76008, 16.740747, 16.734869, 16.739376, 16.75102, 16.765934, 16.780031, 16.788927, 16.788082, 16.774078, 16.744177, 16.697437, 16.634933, 16.557247, 16.464962, 16.358574, 16.240635, 16.1149, 15.989548, 15.875354, 15.779127, 15.701962, 15.645007, 15.608356, 15.5916195, 15.59384, 15.613831, 15.650794, 15.710458, 15.7806015, 15.8631315, 15.955796, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 15.830238, 15.491641, 15.0635195, 14.561173, -999.0, 13.406955, -999.0, -999.0, -999.0, 10.763684, -999.0, 9.235542, -999.0, 7.683046, -999.0, 6.276379, 5.674478, 5.1609716, -999.0, -999.0, -999.0, -999.0, -999.0, 4.06311, 4.194539, 4.400801, 4.667616, 4.979654, 5.320323, 5.6734, 6.0244823, 6.3597894, 6.667956, 6.9391046, 7.164143, 7.336698, 7.451385, 7.50862, 7.5097795, 7.46052, 7.3691, 7.24431, 7.09711, 6.939121, 6.7835712, 6.6441417, 6.532995, 6.462116, 6.442012, 6.480674, 6.585284, 6.757529, 6.9987035, 7.304224, 7.6681056, 8.082257, 8.536109, 9.018083, 9.514665, 10.011977, 10.496422, 10.954472, 11.376621, 11.755019, 12.083075, 12.3567505, 12.573102, 12.733041, 12.838333, 12.894868, 12.909688, 12.889849, 12.842849, 12.776521, 12.69887, 12.617523, 12.5380945, 12.465585, 12.402407, 12.3497305, 12.30869, 12.279824, 12.262998, 12.255942, 12.255769, 12.257389, 12.254547, 12.243479, 12.221148, 12.184036, 12.128487, 12.051086, 11.949568, 11.821892, 11.667791, 11.487933, 11.284559, 11.061706, 10.823224, 10.573377, 10.316792, 10.059659, 9.808616, 9.5700445, 9.350077, 9.153676, 8.983758, 8.843477, 8.735838, 8.663685, 8.627828, 8.6277275, 8.661301, 8.724499, 8.814502, 8.930693, 9.071933, 9.23383, 9.411251, 9.601955, 9.80587, 10.021869, 10.248179, 10.483725, 10.729442, 10.986574, 11.25352, -999.0, 11.803135, 12.078488, 12.348536, 12.607275, 12.848318, 13.064964, 13.250305, 13.398147, 13.503225, 13.560313, 13.565753, 13.516348, 13.412641, 13.256489, 13.051298, 12.802145, 12.514192, 12.193769, 11.8480215, 11.487128, 11.121758, 10.761286, 10.414481, 10.088856, 9.79007, 9.523854, 9.294897, 9.107184, 8.960824, 8.854609, 8.787393, 8.757419, 8.761993, 8.796746, 8.857511, 8.9407, 9.042597, 9.157904, 9.280447, 9.404558, 9.525444, 9.639192, 9.744411, 9.839721, 9.92169, 9.986324, 10.031127, 10.054952, 10.057075, 10.037925, 9.997865, 9.936732, 9.854458, 9.752404, -999.0, 9.496612, 9.344318, 9.176495, 8.995711, 8.805137, 8.60958, 8.414505, 8.204439, 8.019089, 7.841333, 7.6745257, 7.5218754, 7.385861, 7.2689147, 7.1737404, 7.10302, 7.057927, 7.0374613, 7.039951, 7.0616283, 7.098178, 7.144473, 7.1951814, 7.2468643, 7.2975755, 7.344108, 7.381164, 7.403814, 7.409518, 7.3964887, 7.364552, 7.3145933, -999.0, 7.165999, -999.0, -999.0, 6.850593, 6.733804, 6.6156664, 6.501047, 6.3962107, 6.304162, 6.2217636, 6.145775, 6.075413, 6.0104876, 5.949915, 5.8920546, 5.8355136, 5.779243, 5.721448, 5.65795, 5.5845275, 5.5001116, -999.0, 5.2996635, 5.1839995, 5.0588517, 4.9264474, 4.789438, 4.6516933, 4.517608, 4.393328, 4.2863, 4.2038875, 4.153267, 4.140489, 4.16746, 4.235016, 4.34304, 4.490828, 4.6755, 4.891593, 5.132446, 5.388615, 5.650132, 5.906588, 6.1474943, 6.364106, 6.549224, 6.696917, 6.8035913, 6.866812, 6.8881965, 6.8706865, 6.819369, 6.7407694, 6.6436777, 6.5400367, 6.441803, 6.3602166, 6.3060565, 6.2876086, 6.311881, 6.3835096, 6.504667, 6.6759424, 6.8945627, 7.1565065, 7.453483, 7.7757087, 8.112871, 8.372132, 8.704905, 9.023088, 9.315897, 9.573669, 9.787297, 9.950791, 10.0694, 10.119571, 10.116306, 10.061814, 9.962386, 9.824926, 9.657446, 9.469189, 9.27088, 9.074869, 8.892679, 8.732511, 8.602643, 8.510145, 8.461601, 8.462483, 8.51594, 8.623961, 8.783092, 8.989883, 9.238638, 9.522792, 9.834677, 10.165432, 10.505937, 10.846582, 11.177736, 11.490935, 11.777502, 12.030085, 12.242328, 12.4096155, 12.530233, 12.602539, 12.627126, 12.604732, 12.538113, 12.43091, 12.2885, 12.1178255, 11.925311, 11.716919, 11.498801, 11.276914, 11.057002, 10.843121, 10.638433, 10.446206, 10.269213, 10.109647, 9.967774, 9.843655, 9.736433, 9.644819, 9.566887, 9.4999485, 9.440964, 9.386004, 9.33109, 9.27218, 9.205265, 9.126745, 9.033128, 8.920324, 8.783943, 8.620317, 8.428599, 8.208202, 7.9594193, 7.6835194, 7.384099, 7.06616, 6.7303658, 6.3722486, 5.9902925, 5.5994377, 5.218305, 4.855957, 4.5157084, 4.2005863, 3.910527, 3.6464698, 3.4132044, 3.2159138, 3.055549, 2.9310188, 2.841369, 2.7836435, 2.75453, 2.7489448, -999.0, 2.7872055, 2.8249197, 2.8634555, 2.9029133, 2.9395652, 2.9702408, 2.9921033, 3.005042, 3.0095968, 3.0059624, 2.994162, 2.972919, 2.9392445, 2.891077, 2.8285756, 2.7520056, 2.660155, 2.5512917, 2.4232626, 2.2734056, 2.0995662, 1.9024669, 1.6824015, 1.441902, 1.1841767, -999.0, 0.63853556, 0.3637566, 0.09647444, -0.15641405, -0.38795108, -0.5909703, -0.7600106, -0.890175, -0.97662807, -1.01705, -1.0101207, -0.9613586, -0.87710196, -0.76489896, -0.6327041, -0.48489583, -0.32338756, -0.15270059, 0.019395135, 0.18563277, 0.34190002, 0.48409772, 0.60925287, 0.7157606, 0.80289614, 0.8725223, 0.9263592, -999.0, 1.0000358, 1.0275633, 1.0546542, 1.0854512, 1.1235855, 1.1722534, 1.2328446, 1.3074023, 1.3974882, 1.504467, 1.6262848, 1.7580029, 1.8949579, 2.0310388, 2.1601083, 2.2758482, 2.371711, 2.4411929, 2.4777224, 2.4752574, 2.4295154, 2.3362062, 2.1953936, 2.0068905, 1.7740242, 1.5015954, 1.1959012, 0.86581, 0.5202597, 0.169189, -0.1770718, -0.50997317, -0.8207258, -1.1025487, -1.3505564, -1.560907, -1.7351162, -1.8749697, -1.9884645, -2.084039, -2.1707888, -2.2591686, -2.361335, -2.4899533, -2.6550815, -2.8600805, -3.1100771, -3.4117026, -3.7713256, -4.186954, -4.6501255, -5.1537075, -5.688008, -6.242703, -6.8050547, -7.361426, -7.898653, -8.403817, -8.866988, -9.32204, -9.680694, -999.0, -10.226825, -10.407123, -10.520667, -10.567838, -10.552187, -10.478313, -10.354212, -10.187676, -9.986704, -9.759303, -9.514472, -9.261564, -9.010994, -8.773957, -8.560923, -8.379544, -8.237562, -8.140819, -8.094403, -8.1006565, -8.159524, -8.270127, -8.429123, -8.632764, -8.875602, -9.151952, -9.456089, -9.782017, -10.122572, -10.469589, -10.815743, -11.155482, -11.483244, -11.793193, -12.079586, -12.337675, -12.563404, -12.752852, -12.9028635, -13.010848, -13.076818, -13.101463, -13.08731, -13.037999, -12.957322, -12.849817, -12.72078, -12.577755, -12.428639, -12.281308, -12.143522, -12.020857, -11.916857, -11.835145, -11.778294, -11.748358, -11.744126, -11.763486, -11.802907, -11.857436, -11.921706, -11.989485, -12.054394, -12.111327, -12.155616, -12.1865635, -12.205612, -12.2146225, -12.21711, -12.216847, -12.219405, -12.230838, -12.259032, -12.312684, -12.399532, -12.526204, -12.697945, -12.915621, -13.179863, -13.488043, -13.836526, -14.218914, -14.626545, -15.050071, -15.478297, -15.899731, -16.302715, -16.675694, -17.009481, -17.321741, -17.548695, -17.716936, -17.823074, -17.866465, -17.846882, -17.767078, -17.630638, -17.44371, -17.214016, -16.949104, -16.656681, -16.34443, -16.019205, -15.687653, -15.354351, -15.023059, -14.69679, -14.377335, -14.065598, -13.760535, -13.461048, -13.167297, -12.879807, -12.600774, -12.33356, -12.080863, -11.845066, -11.628864, -11.436334, -11.271886, -11.140477, -11.04738, -10.996599, -10.990254, -11.029984, -11.114132, -11.240492, -11.403897, -11.598198, -11.817571, -12.055676, -12.304961, -12.55626, -12.800656, -13.032562, -13.247025, -13.441784, -13.616557, -13.770804, -13.905585, -14.022828, -14.129041, -14.2322855, -14.342097, -14.467817, -14.610801, -14.765467, -14.930704, -15.113227, -15.320039, -15.554802, -15.820489, -16.113817, -16.426008, -16.74965, -17.077168, -17.40058, -17.71233, -18.004827, -18.271519, -18.506641, -18.705435, -18.865349, -18.98371, -19.060167, -19.09466, -19.090067, -19.050497, -18.98056, -18.886005, -18.772772, -18.646803, -18.513962, -18.37833, -18.24366, -18.113209, -17.989618, -17.875269, -17.771479, -17.679361, -17.598242, -17.527025, -17.463648, -17.405567, -17.351175, -17.299835, -17.251001, -17.204771, -17.161158, -17.120003, -17.081244, -17.04251, -17.012539, -16.988773, -16.972086, -16.963467, -16.963789, -16.973791, -16.993193, -17.021343, -17.05728, -17.099644, -17.147055, -17.197891, -17.250246, -17.301414, -17.348736, -17.391003, -999.0, -17.456854, -17.476282, -17.48422, -17.481329, -17.468716, -17.448774, -17.424522, -17.399736, -999.0, -17.36567, -17.363495, -17.375603, -17.406008, -17.458986, -17.539083, -17.650707, -17.794832, -17.96779, -18.164312, -18.375462, -18.592718, -18.813543, -19.037186, -19.25722, -19.462269, -19.641415, -19.784266, -19.880863, -19.923597, -19.9053, -19.818512, -19.65671, -19.421112, -999.0, -18.96052, -18.60669, -18.238676, -17.872223, -17.514378, -17.17218, -16.855268, -16.573662, -16.336275, -16.151138, -16.023418, -15.953389, -15.94031, -15.979279, -16.06388, -16.183647, -16.326235, -16.48267, -16.647173, -16.812672, -16.969858, -17.109783, -17.227242, -17.318289, -17.380047, -17.411253, -17.412086, -17.385954, -17.33657, -17.268423, -999.0, -17.094385, -16.997414, -16.901562, -16.814999, -16.744595, -16.69271, -16.661264, -16.652739, -16.66948, -16.712927, -16.78284, -16.878183, -16.994263, -17.125517, -17.26492, -17.405024, -17.541927, -17.674751, -17.801685, -17.931122, -18.036137, -18.12499, -18.19348, -18.239895, -18.26383, -18.265776, -18.248339, -18.214415, -999.0, -18.111633, -18.048216, -17.97936, -17.908945, -17.84181, -17.781075, -17.727125, -17.680887, -17.643934, -999.0, -17.601458, -17.593918, -17.593445, -17.598152, -17.606672, -17.61819, -17.63129, -17.641844, -17.64518, -17.64027, -17.628872, -17.611263, -17.58633, -999.0, -17.514387, -17.471552, -17.427752, -17.386377, -17.350826, -17.32468, -17.311428, -17.31396, -17.335226, -17.378092, -17.445105, -17.537037, -17.652617, -17.790985, -17.951067, -18.13159, -18.328793, -18.537981, -18.752838, -18.965214, -19.166418, -19.347906, -19.502413, -19.629217, -19.728922, -19.801472, -19.846851, -19.864088, -19.850868, -19.805191, -19.726847, -19.615643, -19.47406, -19.306707, -999.0, -18.943256, -999.0, -18.612106, -18.461542, -18.321482, -18.193102, -18.08198, -17.995762, -17.936756, -17.90057, -999.0, -17.886011, -17.90502, -17.935728, -17.971497, -18.007523, -18.040607, -18.067806, -999.0, -18.098625, -18.099579, -18.08932, -18.068344, -18.038935, -999.0, -17.969511, -17.940989, -17.925146, -17.928274, -17.952524, -17.997702, -18.064627, -18.154392, -18.280613, -18.42014, -18.582588, -18.764256, -18.960787, -19.168633, -19.383627, -19.598505, -19.802137, -19.984835, -20.144522, -20.280416, -20.392487, -20.481714, -20.547884, -20.5898, -20.607164, -20.602392, -20.578083, -20.537447, -20.484158, -20.422033, -20.355206, -999.0, -20.225508, -20.171923, -20.129786, -20.100784, -20.084112, -20.077015, -20.077791, -999.0, -20.099924, -20.118618, -20.140465, -20.165157, -20.192759, -20.222233, -20.251131, -999.0, -999.0, -20.296572, -20.294146, -20.27897, -20.249662, -20.20251, -20.13414, -20.046797, -19.94524, -19.83487, -19.721834, -19.609844, -19.497435, -19.383484, -19.271412, -19.165674, -19.071083, -18.993397, -18.938007, -999.0, -18.907877, -18.936007, -18.992363, -999.0, -999.0, -19.305374, -19.446833, -19.60048, -19.759085, -19.915144, -20.062775, -20.196594, -20.312853, -20.409796, -20.48592, -20.540583, -20.572678, -20.580257, -20.561516, -20.518261, -20.454535, -20.373789, -20.27958, -20.175783, -20.066376, -19.95514, -19.844292, -19.735481, -999.0, -19.535168, -19.449432, -19.375267, -19.31382, -19.26615, -19.233212, -19.215801, -19.214334, -19.228273, -19.25602, -19.29654, -19.351576, -19.423677, -19.515207, -19.62802, -19.760057, -19.904451, -20.055882, -20.212505, -20.372736, -20.53439, -20.695019, -20.850048, -20.993273, -21.132074, -21.240238, -21.330057, -21.399704, -21.447159, -21.470425, -21.467678, -999.0, -21.38603, -21.310863, -21.214989, -21.100807, -20.974575, -20.843718, -20.712227, -20.581396, -20.453505, -20.331005, -20.215712, -20.108389, -999.0, -19.966, -19.889627, -999.0, -19.791473, -19.760801, -19.73858, -19.724508, -19.717224, -19.715328, -19.717852, -19.726105, -19.741926, -19.766174, -19.799215, -19.840805, -19.889248, -19.9432, -999.0, -20.06046, -20.118317, -20.170746, -20.214607, -20.246367, -20.261171, -20.252373, -20.212963, -20.14055, -20.03462, -19.900248, -19.746351, -19.57698, -19.390491, -19.186983, -18.972073, -18.751698, -999.0, -18.315928, -18.112612, -17.92774, -17.766743, -17.631554, -17.524336, -17.447449, -17.402784, -17.389225, -17.403202, -17.441748, -17.50219, -17.582043, -999.0, -17.789288, -17.908825, -18.031368, -18.151825, -18.266062, -18.370455, -18.463224, -18.54239, -18.604784, -18.64718, -18.669163, -18.672983, -18.660213, -18.632635, -18.592701, -18.544933, -18.49405, -18.442198, -18.390173, -18.340248, -18.296179, -18.261541, -18.2382, -18.227541, -18.228594, -18.239107, -18.257957, -999.0, -18.32222, -18.370815, -18.432922, -999.0, -18.553068, -18.635736, -18.722338, -18.811527, -18.902275, -18.99384, -19.085236, -19.175241, -19.262505, -19.345013, -19.420492, -19.486485, -19.540495, -19.58168, -19.610342, -19.62693, -19.632635, -19.628572, -19.615513, -19.594193, -19.56537, -19.5298, -19.48854, -19.442942, -19.394192, -19.343517, -999.0, -19.242062, -19.195345, -19.154757, -19.123089, -19.101595, -19.089235, -19.085506, -19.091253, -19.10742, -19.134043, -19.170612, -19.21547, -19.266052, -19.32155, -19.384188, -19.45555, -19.532322, -19.609951, -999.0, -19.759762, -19.830141, -19.89718, -19.961, -20.021454, -20.077953, -20.127625, -20.16668, -20.194534, -999.0, -20.228262, -20.236555, -20.239178, -20.235928, -20.226631, -20.213234, -20.199497, -20.188007, -20.179155, -20.173355, -20.17103, -20.1725, -20.178066, -20.187931, -20.201895, -20.219051, -20.238586, -20.259577, -20.28101, -20.30123, -20.318157, -20.329523, -20.333035, -20.326962, -20.31169, -999.0, -20.272934, -20.238428, -20.19915, -20.157549, -20.115688, -20.073303, -20.029467, -19.986044, -19.947407, -19.917072, -19.894758, -19.88535, -19.884527, -19.890055, -19.900646, -19.915102, -19.931087, -19.945293, -19.955055, -19.959684, -999.0, -19.95113, -19.935968, -19.911499, -19.875875, -19.828169, -19.771091, -19.707918, -19.644049, -19.585594, -19.536364, -19.498486, -19.474342, -19.46575, -19.474337, -19.500978, -999.0, -19.614717, -19.706997, -19.821667, -19.95076, -20.08758, -20.22757, -20.36619, -20.500183, -20.62681, -20.742096, -20.841536, -20.921768, -20.982128, -21.021942, -21.041624, -21.04208, -21.02501, -20.992651, -999.0, -20.888893, -20.819508, -20.739538, -20.650345, -999.0, -20.512474, -20.428644, -20.356386, -20.298897, -20.255583, -20.223068, -20.199226, -20.182701, -20.17202, -20.165741, -20.162447, -999.0, -20.15546, -20.146132, -20.129082, -20.102392, -20.067146, -20.024632, -19.975786, -19.921364, -19.860693, -19.792284, -19.715994, -19.633959, -999.0, -19.465168, -19.3843, -19.301949, -19.210533, -19.108866, -19.00226, -18.894503, -18.785902, -18.676636, -999.0, -18.443455, -18.312122, -18.168606, -18.013227, -17.851185, -17.686909, -999.0, -17.435602, -17.26483, -17.094818, -16.928408, -16.767145, -16.61284, -16.468739, -16.338245, -16.222887, -16.119644, -16.01657, -15.930396, -15.849642, -999.0, -15.705038, -999.0, -15.582276, -15.525793, -15.47006, -15.413026, -15.35306, -15.288148, -15.2158785, -15.134814, -15.046466, -14.956524, -14.869329, -14.782028, -14.690796, -14.594123, -14.490898, -14.379956, -14.261931, -14.139151, -14.015248, -13.893575, -13.769115, -13.633009, -13.478004, -999.0, -13.09879, -12.884189, -999.0, -12.431001, -12.182329, -11.918524, -11.643916, -11.359011, -11.062908, -10.757348, -10.451985, -10.157421, -9.877288, -9.61223, -9.362142, -999.0, -8.898352, -8.68538, -8.487314, -8.304073, -8.13556, -7.9817786, -999.0, -7.7124534, -7.5891395, -999.0, -7.3514915, -7.2431955, -7.144537, -7.0564985, -6.9801745, -6.9161515, -6.864949, -6.826476, -6.8007092, -6.787776, -6.787874, -6.800348, -999.0, -6.8542314, -6.890004, -6.9272904, -6.962273, -6.9905124, -7.0062213, -7.0031724, -6.977722, -6.929944, -6.858412, -6.760199, -999.0, -6.4772677, -6.2973537, -6.096622, -5.8804626, -5.6544566, -5.424839, -5.1975946, -4.9770265, -4.76706, -4.5731926, -999.0, -4.3275976, -4.2045956, -4.122038, -4.080083, -4.07178, -4.0918164, -4.1357055, -4.1981497, -4.2726707, -4.352964, -4.4440365, -4.527584, -4.608356, -4.6813803, -4.74204, -4.7873645, -4.8145747, -4.8243556, -999.0, -4.8013525, -4.776183, -4.747621, -4.7197003, -4.696587, -4.682072, -999.0, -4.69277, -4.723249, -4.773038, -4.842379, -4.931425, -5.0384517, -5.1612616, -5.296131, -999.0, -5.58422, -5.7290854, -5.8694763, -6.003137, -6.127578, -6.2402587, -6.338899, -6.4234223, -6.495561, -6.5570345, -6.6099215, -6.6561365, -6.696318, -6.730893, -6.7601867, -6.7843146, -6.8033614, -6.8173428, -6.8262787, -6.830328, -6.8295856, -6.8244348, -6.8155026, -6.804404, -6.7936244, -6.7853255, -6.780819, -6.781156, -6.785688, -6.7933183, -6.8027816, -6.812565, -6.8212814, -6.8276844, -6.830619, -999.0, -6.820259, -6.802477, -6.7720985, -6.7269917, -6.6664653, -6.5909653, -6.5034547, -6.4060416, -6.2975316, -6.1765037, -999.0, -5.9813433, -5.8526535, -5.7293916, -5.613387, -5.505716, -5.405935, -5.3143435, -5.2327104, -5.162637, -5.104993, -5.060586, -5.03061, -5.016484, -5.0194793, -5.0406933, -5.082003, -5.1450853, -5.230792, -5.335617, -5.454194, -5.58576, -5.7349067, -5.904629, -6.094342, -6.30354, -6.531896, -6.778836, -7.044228, -7.3279324, -7.6278176, -7.9405627, -8.265648, -8.608929, -999.0, -9.36291, -9.755468, -10.14537, -10.526029, -10.889829, -11.2297535, -11.539024, -11.840271, -12.078094, -12.282896, -12.457155, -12.599644, -12.703436, -12.762778, -12.778428, -12.752162, -12.686699, -12.585863, -12.452301, -12.288123, -12.097113, -11.886459, -11.662682, -11.427259, -11.180727, -10.928761, -10.67996, -10.438332, -10.2006645, -9.965222, -9.737522, -9.524222, -9.328136, -9.150125, -8.99095, -999.0, -8.725982, -8.618005, -8.525017, -8.44858, -8.391587, -8.355891, -999.0, -8.348772, -8.373573, -8.41341, -8.467287, -8.53442, -8.611946, -8.695321, -8.780053, -8.861844, -8.93667, -9.003251, -9.060758, -9.108318, -9.145484, -9.172311, -9.190211, -9.200892, -9.207751, -9.214551, -9.224628, -9.241236, -9.266657, -9.301597, -9.3466015, -9.400661, -9.462656, -9.531016, -9.603849, -9.679076, -9.754651, -9.82917, -9.902816, -9.975879, -10.049146, -10.123329, -10.1982, -10.273349, -10.35001, -10.430969, -10.518069, -10.611091, -10.709708, -10.814847, -10.927828, -11.05075, -11.18663, -11.337937, -11.505792, -11.69152, -11.895909, -12.119521, -12.361881, -12.621832, -12.898835, -13.191833, -13.499301, -13.815961, -14.136339, -14.454541, -14.763855, -15.056921, -15.324907, -15.557979, -15.746369, -15.880657, -15.958325, -15.976939, -15.929524, -15.817971, -15.643422, -15.415201, -15.142376, -14.838396, -14.517806, -14.195332, -13.886044, -13.603504, -13.359264, -13.165579, -13.031784, -12.967302, -12.973045, -999.0, -13.178738, -13.355868, -13.56958, -13.817067, -14.09363, -14.3869, -14.683034, -14.965632, -15.2171335, -15.424822, -15.581008, -15.6779785, -15.711554, -15.679371, -15.5877285, -15.445461, -999.0, -15.045072, -14.80586, -14.552399, -14.2924595, -14.030269, -13.769272, -13.51211, -13.261003, -13.018526, -12.786543, -12.564026, -12.342972, -12.115011, -999.0, -11.619528, -999.0, -11.050749, -10.739253, -10.419827, -10.099847, -9.781714, -9.468653, -9.173927, -999.0, -8.703051, -8.540118, -8.429359, -999.0, -8.373356, -8.434762, -8.561583, -8.751923, -999.0, -9.290931, -9.626263, -9.995671, -10.384138, -999.0, -999.0, -11.333714, -11.667984, -11.953772, -12.175573, -12.322371, -12.388974, -12.372951, -12.281172, -12.121151, -999.0, -11.776373, -11.494106, -999.0, -10.874021, -10.576417, -10.319773, -10.123414, -999.0, -9.956864, -9.993204, -10.122681, -10.317983, -999.0, -10.902416, -11.266827, -11.665499, -12.089538, -12.520036, -12.918411, -13.248159, -13.496879, -999.0, -13.732524, -13.717164, -13.611051, -13.40936, -13.109256, -12.718743, -12.25142, -999.0, -11.491722, -11.0119705, -10.584005, -999.0, -9.935349, -9.709202, -9.546923, -9.45807, -9.450769, -9.527893, -999.0, -9.794787, -10.043591, -999.0, -10.636682, -10.976788, -999.0, -11.692868, -12.040201, -12.366963, -12.66193, -999.0, -13.009509, -13.160421, -13.244171, -999.0, -999.0, -13.077154, -12.883168, -12.631506, -12.333107, -12.0012245, -11.648836, -11.287883, -10.928963, -999.0, -10.234669, -9.912012, -999.0, -999.0, -9.184124, -999.0, -8.976537, -8.973133, -9.04291, -9.188912, -9.4033165, -9.663691, -9.948946, -10.2451935, -999.0, -10.832324, -11.121088, -999.0, -11.69126, -11.966173, -12.214472, -12.418441, -12.568736, -12.658518, -12.686184, -999.0, -999.0, -999.0, -12.363834, -12.178098, -11.962051, -11.726248, -11.490857, -11.27539, -11.088758, -10.9363365, -10.819775, -999.0, -999.0, -10.682721, -10.699712, -10.761708, -10.866205, -11.009185, -11.182639, -11.377596, -999.0, -999.0, -999.0, -12.068822, -12.225661, -999.0, -12.433747, -999.0, -12.475001, -12.425571, -12.319211, -999.0, -12.050924, -999.0, -11.684613, -11.44519, -11.213091, -10.993175, -10.782688, -999.0, -10.396127, -999.0, -10.096927, -9.995016, -999.0, -9.885937, -9.8709755, -999.0, -9.913523, -9.966591, -10.036206, -10.118362, -10.208706, -10.302815, -10.396444, -10.486707, -10.5743885, -10.660475, -10.744084, -10.823872, -10.899955, -10.973621, -11.046014, -11.117879, -999.0, -11.224434, -11.291665, -11.35485, -999.0, -11.483325, -11.554208, -11.631233, -999.0, -11.795801, -11.877379, -11.956954, -999.0, -12.098643, -12.148392, -12.181288, -12.199647, -12.204364, -12.194965, -12.172063, -12.139422, -12.101768, -12.06663, -12.042525, -12.035667, -999.0, -12.091885, -12.170672, -12.286495, -999.0, -12.660009, -12.911802, -13.184475, -13.463731, -999.0, -999.0, -14.266477, -14.504914, -14.728567, -14.942063, -15.137662, -999.0, -15.355649, -15.431947, -15.446337, -15.397989, -999.0, -999.0, -14.938821, -14.721031, -999.0, -14.235892, -13.975337, -13.710116, -13.446248, -13.189875, -12.947239, -12.724971, -12.529686, -12.366536, -12.239674, -12.151171, -12.097094, -12.086604, -999.0, -12.1782465, -12.278157, -12.409489, -12.564579, -12.732707, -12.9083605, -13.09533, -13.294785, -13.493311, -13.674788, -999.0, -13.971084, -14.084728, -14.168975, -14.218296, -14.22849, -14.196771, -14.128745, -999.0, -13.977659, -13.851347, -13.707966, -13.55325, -13.394534, -13.240126, -13.099484, -12.980475, -12.886474, -12.819954, -12.782383, -12.7747345, -12.796238, -999.0, -12.917148, -13.011056, -999.0, -13.246128, -13.374362, -13.501145, -13.620557, -13.729409, -13.828409, -13.916905, -13.988867, -14.038082, -14.065638, -14.076093, -14.073239, -14.06003, -14.037968, -999.0, -13.9602375, -13.903824, -999.0, -13.766365, -13.693112, -13.623276, -13.562669, -13.516292, -999.0, -999.0, -999.0, -999.0, -999.0, -13.545186, -999.0, -13.674018, -13.759151, -999.0, -13.960283, -14.071588, -14.18631, -14.301378, -999.0, -999.0, -14.616299, -14.704093, -999.0, -999.0, -14.888149, -14.915398, -14.92725, -14.9258995, -999.0, -14.891624, -14.8580065, -999.0, -14.758839, -14.703983, -14.648848, -14.59179, -14.532341, -14.471705, -14.411705, -999.0, -14.306406, -14.259393, -14.207142, -14.147706, -14.084812, -14.015074, -999.0, -13.889249, -999.0, -13.770175, -13.720197, -999.0, -13.670639, -13.677897, -13.709175, -13.767018, -999.0, -13.906334, -999.0, -14.169048, -14.323189, -999.0, -14.654174, -14.81626, -14.967989, -15.10706, -15.20555, -15.318874, -999.0, -15.49967, -15.559592, -15.594349, -15.60227, -15.583775, -15.545073, -15.492985, -15.4323635, -15.367086, -999.0, -15.220314, -15.13792, -15.059438, -14.994027, -14.9467745, -14.921563, -14.917101, -14.928166, -999.0, -14.986328, -15.0310545, -15.084045, -15.143968, -15.210612, -999.0, -15.360112, -15.43329, -999.0, -15.555128, -15.604089, -15.647952, -999.0, -15.7309, -15.768772, -15.800433, -999.0, -15.8215275, -999.0, -999.0, -999.0, -999.0, -999.0, -15.544603, -15.465394, -15.385542, -15.305653, -999.0, -15.153086, -15.086131, -999.0, -14.9875345, -14.958784, -14.942102, -999.0, -14.953331, -14.986941, -999.0, -15.093445, -15.154714, -999.0, -15.239224, -15.287743, -15.329879, -15.363875, -999.0, -15.400854, -15.403471, -15.396865, -999.0, -15.368034, -15.349671, -15.32943, -15.308239, -999.0, -999.0, -15.255352, -999.0, -15.251393, -15.259634, -15.277328, -15.308644, -15.354358, -15.410963, -15.475371, -15.545249, -15.618325, -15.692526, -15.765753, -999.0, -15.894248, -15.945036, -999.0, -15.98684, -15.974842, -15.934152, -15.864676, -15.768771, -999.0, -15.500996, -15.33183, -15.14564, -14.948629, -14.745033, -14.537597, -14.322975, -14.093758, -999.0, -999.0, -13.371417, -13.154778, -12.959954, -999.0, -12.720039, -999.0, -999.0, -999.0, -12.4434805, -999.0, -999.0, -12.560252, -12.654722, -12.766284, -999.0, -999.0, -999.0, -13.352095, -13.559646, -13.789794, -14.023224, -14.240933, -14.441668, -14.630103, -14.804924, -14.962081, -999.0, -999.0, -15.337973, -15.443835, -999.0, -15.642084, -15.742652, -15.850842, -999.0, -999.0, -16.18129, -16.342485, -999.0, -999.0, -16.871878, -999.0, -17.230997, -17.41955, -999.0, -17.702478, -17.874182, -18.013002, -18.11505, -999.0, -18.23561, -18.2606, -999.0, -18.245811, -999.0, -999.0, -18.117353, -18.052069, -17.982388, -17.906261, -999.0, -17.748493, -17.674093, -17.600216, -999.0, -999.0, -999.0, -17.322308, -17.232582, -17.134333, -17.028273, -16.916546, -999.0, -16.695297, -999.0, -16.51675, -16.444752, -16.385185, -999.0, -999.0, -16.199734, -16.156553, -16.13165, -16.128536, -16.148651, -16.194677, -16.26968, -999.0, -999.0, -999.0, -16.747736, -999.0, -17.109283, -17.302067, -999.0, -17.692728, -17.877111, -999.0, -999.0, -18.24584, -999.0, -18.40488, -18.430054, -999.0, -18.36857, -18.278137, -999.0, -17.954145, -999.0, -999.0, -17.294313, -16.9986, -16.712627, -16.428701, -16.139143, -15.849597, -999.0, -999.0, -999.0, -999.0, -14.794653, -14.669279, -14.594743, -14.562902, -14.5681505, -14.608989, -999.0, -14.797221, -14.947511, -15.126279, -15.314996, -15.500959, -15.679006, -15.8424, -999.0, -16.093348, -16.166655, -16.198328, -999.0, -16.13505, -999.0, -16.006231, -15.904849, -15.803966, -15.709526, -15.62924, -15.572549, -15.549074, -15.563518, -15.617325, -15.710249, -15.836946, -999.0, -16.174633, -999.0, -999.0, -16.773222, -999.0, -17.110641, -17.249624, -17.362394, -17.44425, -17.492334, -17.504248, -17.478613, -999.0, -17.30932, -17.159302, -16.96116, -16.719868, -999.0, -999.0, -16.024221, -15.775211, -15.546203, -15.324024, -15.106731, -14.896192, -14.698991, -14.529557, -14.39854, -999.0, -14.270832, -14.229372, -14.221232, -14.243561, -999.0, -999.0, -999.0, -14.480049, -14.538812, -14.581446, -14.602318, -999.0, -14.565381, -14.502718, -14.404478, -14.281536, -14.152042, -14.020212, -13.875152, -13.712273, -999.0, -13.4587965, -13.29472, -13.131178, -12.96628, -12.805447, -12.654745, -12.515418, -999.0, -999.0, -999.0, -999.0, -12.009597, -999.0, -11.83943, -11.761539, -11.686125, -999.0, -11.55783, -11.509195, -11.469479, -999.0, -999.0, -11.401979, -11.381193, -11.357272, -11.325636, -11.282988, -11.227832, -11.164524, -11.097434, -11.024515, -10.941442, -999.0, -999.0, -999.0, -10.622457, -10.551929, -10.502936, -10.480971, -10.491431, -999.0, -999.0, -999.0, -999.0, -10.91111, -11.07052, -999.0, -11.428572, -11.6136055, -11.7922125, -11.9576645, -999.0, -12.230478, -12.335641, -999.0, -12.474185, -12.502258, -12.499381, -12.465238, -12.405284, -12.324901, -12.226771, -12.112908, -11.985782, -11.848723, -999.0, -11.575316, -11.460694, -11.369074, -11.304882, -11.272543, -11.275529, -999.0, -999.0, -999.0, -11.553681, -11.684299, -11.827317, -11.98564, -12.157935, -12.330796, -999.0, -12.633654, -12.7601595, -12.874045, -12.946215, -12.984662, -999.0, -12.974415, -12.929978, -12.859374, -999.0, -12.626113, -12.465552, -999.0, -12.209533, -999.0, -11.893681, -11.759021, -11.644054, -11.551487, -999.0, -11.436938, -999.0, -11.4030905, -999.0, -11.419926, -11.441175, -999.0, -999.0, -999.0, -11.562791, -11.57467, -11.569385, -11.546602, -999.0, -11.494474, -11.455041, -11.412856, -999.0, -11.318616, -999.0, -11.203698, -11.142022, -999.0, -999.0, -11.008125, -10.972911, -10.950051, -10.939155, -999.0, -999.0, -10.947956, -999.0, -999.0, -10.950494, -999.0, -999.0, -10.894803, -10.848661, -999.0, -999.0, -10.63183, -10.537806, -10.437869, -10.334725, -10.22722, -10.1135025, -999.0, -9.879438, -9.7696295, -999.0, -999.0, -999.0, -9.470938, -999.0, -9.4184265, -999.0, -9.410868, -9.415718, -999.0, -9.439163, -999.0, -9.467724, -9.478485, -9.485579, -999.0, -9.489793, -999.0, -999.0, -999.0, -9.490987, -9.48878, -9.4826975, -9.471493, -999.0, -999.0, -999.0, -9.391624, -9.374804, -999.0, -9.357329, -999.0, -9.359416, -9.362866, -9.364123, -999.0, -9.358183, -9.350674, -999.0, -9.330231, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -8.970845, -8.866695, -999.0, -8.719827, -999.0, -999.0, -8.5195465, -8.467259, -8.419153, -999.0, -8.361702, -999.0, -8.348788, -8.355681, -999.0, -999.0, -8.448452, -999.0, -8.578495, -8.65761, -999.0, -8.83344, -8.92641, -999.0, -9.065556, -9.150914, -999.0, -9.285136, -9.33598, -999.0, -999.0, -999.0, -9.470461, -999.0, -9.48977, -9.488469, -9.484405, -9.486722, -9.504685, -999.0, -999.0, -999.0, -9.727095, -999.0, -9.779999, -999.0, -9.047951, -999.0, -999.0, -999.0, -999.0, -999.0, -1.0990872, -0.2784979, 0.17485751, -999.0, -999.0, -999.0, -999.0, 0.21400143, 0.053198356, -999.0}
wspd =
  {2.7, -999.0, -999.0, 12.606418, 14.382931, -999.0, -999.0, -999.0, 16.388268, 16.539232, 16.747799, 17.032719, 17.343359, 17.652035, 17.94358, 18.199255, 18.412317, 18.578987, 18.698565, 18.77377, 18.807709, 18.804836, 18.769907, 18.708559, 18.626656, 18.53076, 18.427784, 18.323921, 18.224546, 18.134663, 18.057087, 17.99453, 17.947342, 17.915255, 17.896759, 17.889128, 17.889187, 17.892717, 17.895432, 17.893248, 17.881977, 17.858406, 17.819939, 17.765436, 17.695465, 17.61036, 17.510826, 17.397367, 17.272104, 17.138329, 17.00426, 16.88106, 16.77594, 16.690464, 16.62613, 16.582909, 16.560251, 16.557241, 16.572783, 16.606153, 16.663147, 16.73272, 16.81792, 16.917957, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 17.11896, 16.832174, 16.458178, 16.008446, -999.0, 14.944394, -999.0, -999.0, -999.0, 12.412326, -999.0, 10.926929, -999.0, 9.432717, -999.0, 8.115949, 7.572457, 7.124663, -999.0, -999.0, -999.0, -999.0, -999.0, 6.328115, 6.4575076, 6.643886, 6.87519, 7.138954, 7.4220076, 7.7107844, 7.993281, 8.257524, 8.493843, 8.694002, 8.850623, 8.959319, 9.01636, 9.023062, 8.981837, 8.899076, 8.783709, 8.645279, 8.4952, 8.345571, 8.20922, 8.0992155, 8.02632, 8.000603, 8.030643, 8.122378, 8.280509, 8.50389, 8.791239, 9.136456, 9.532389, 9.970289, 10.439373, 10.928168, 11.423968, 11.91357, 12.384517, 12.824217, 13.224135, 13.577441, 13.879042, 14.127004, 14.320602, 14.46328, 14.559116, 14.615139, 14.639509, 14.641186, 14.629913, 14.615151, 14.605461, 14.6089735, 14.631184, 14.676893, 14.748409, 14.846621, 14.971058, 15.119132, 15.287159, 15.469158, 15.658644, 15.848902, 16.051182, 16.222916, 16.378283, 16.511848, 16.617752, 16.691082, 16.73053, 16.73546, 16.707867, 16.65125, 16.570913, 16.474352, 16.369276, 16.264364, 16.168743, 16.09199, 16.043667, 16.031357, 16.060875, 16.1369, 16.261326, 16.435408, 16.656803, 16.921732, 17.222878, 17.551262, 17.900837, 18.2679, 18.646805, 19.02722, 19.39876, 19.75435, 20.087908, 20.395494, 20.676182, 20.929327, 21.15617, 21.358337, 21.538458, 21.699532, 21.843582, -999.0, 22.085732, 22.18594, 22.27262, 22.3435, 22.395643, 22.426058, 22.43156, 22.409998, 22.360619, 22.282335, 22.174639, 22.037476, 21.87359, 21.686916, 21.48269, 21.267529, 21.048157, 20.831352, 20.623936, 20.431927, 20.260763, 20.114267, 19.994898, 19.903336, 19.838013, 19.79671, 19.775728, 19.77093, 19.777256, 19.789413, 19.801752, 19.808464, 19.804853, 19.78794, 19.754688, 19.702082, 19.627405, 19.530647, 19.413803, 19.281351, 19.14041, 18.99487, 18.841074, 18.675407, 18.500595, 18.321186, 18.140348, 17.96071, 17.784565, 17.613375, 17.448734, 17.292526, 17.146664, 17.011887, -999.0, 16.775236, 16.672863, 16.580614, 16.497828, 16.423765, 16.357529, 16.297766, 16.236225, 16.179913, 16.120106, 16.055492, 15.984746, 15.906763, 15.82072, 15.726551, 15.624417, 15.512312, 15.386142, 15.244134, 15.090992, 14.932849, 14.777472, 14.632383, 14.496567, 14.36224, 14.225999, 14.091966, 13.9642315, 13.845502, 13.738248, 13.644199, 13.564743, -999.0, 13.457635, -999.0, -999.0, 13.453732, 13.495647, 13.557731, 13.636308, 13.725221, 13.819203, 13.915563, 14.011363, 14.10074, 14.177034, 14.234382, 14.26749, 14.272039, 14.245008, 14.183981, 14.088044, 13.956923, 13.792649, -999.0, 13.378303, 13.137862, 12.883172, 12.621908, 12.361998, 12.111536, 11.87864, 11.6709795, 11.4958315, 11.359804, 11.26851, 11.226655, 11.23591, 11.296981, 11.407233, 11.562228, 11.75586, 11.979932, 12.225427, 12.4814415, 12.736441, 12.978124, 13.193839, 13.372769, 13.505789, 13.585234, 13.60626, 13.565377, 13.463736, 13.30411, 13.0922165, 12.835754, 12.544509, 12.231174, 11.909079, 11.592568, 11.296196, 11.033129, 10.815907, 10.65535, 10.560246, 10.537162, 10.587913, 10.712478, 10.9067335, 11.164442, 11.476424, 11.741547, 12.115949, 12.511439, 12.915908, 13.317974, 13.706973, 14.075648, 14.452991, 14.767233, 15.05344, 15.311019, 15.540044, 15.740145, 15.911994, 16.056566, 16.174786, 16.26811, 16.336987, 16.381273, 16.400734, 16.395485, 16.366188, 16.314974, 16.24573, 16.163227, 16.07347, 15.982973, 15.898891, 15.828313, 15.778267, 15.754944, 15.762413, 15.80176, 15.872295, 15.970317, 16.091417, 16.230804, 16.383669, 16.54463, 16.707567, 16.867405, 17.019594, 17.160015, 17.285374, 17.392344, 17.47737, 17.536516, 17.56557, 17.561426, 17.52067, 17.442173, 17.325197, 17.17096, 16.982204, 16.762575, 16.517328, 16.25215, 15.9736, 15.688534, 15.403531, 15.125021, 14.858401, 14.60778, 14.376248, 14.164495, 13.972853, 13.800178, 13.644817, 13.504085, 13.374694, 13.253803, 13.139068, 13.028523, 12.921107, 12.81621, 12.714491, 12.617357, 12.526814, 12.445351, 12.375389, 12.3204565, 12.284503, 12.268903, 12.271985, 12.29289, 12.331806, 12.386717, 12.453218, 12.527243, 12.604922, 12.682164, 12.755628, 12.822741, 12.880934, 12.928132, 12.963065, 12.986264, -999.0, 12.999941, 12.989234, 12.968843, 12.939201, 12.901378, 12.857137, 12.8080015, 12.755174, 12.699946, 12.644453, 12.591094, 12.54146, 12.497018, 12.460311, 12.436082, 12.429215, 12.441611, 12.474422, 12.529589, 12.608924, 12.71422, 12.846265, 13.0060215, 13.193278, 13.407447, -999.0, 13.908238, 14.1869, 14.475949, 14.768432, 15.0561, 15.330273, 15.581615, 15.8000965, 15.975118, 16.097208, 16.158484, 16.159706, 16.102608, 15.992157, 15.834015, 15.630214, 15.381505, 15.092475, 14.77572, 14.442995, 14.105111, 13.773333, 13.457236, 13.16515, 12.9049015, 12.681413, 12.49982, -999.0, 12.261929, 12.202328, 12.17746, 12.182212, 12.208977, 12.250559, 12.299826, 12.349158, 12.391379, 12.419362, 12.428296, 12.415437, 12.378344, 12.317536, 12.233188, 12.127676, 12.0033455, 11.863285, 11.711335, 11.552028, 11.391208, 11.235127, 11.089377, 10.960499, 10.853843, 10.774614, 10.727498, 10.7152195, 10.739304, 10.797642, 10.886568, 10.999725, 11.129268, 11.266926, 11.404313, 11.533396, 11.647737, 11.740952, 11.809089, 11.848754, 11.860406, 11.84646, 11.810208, 11.757161, 11.693541, 11.626804, 11.565069, 11.517658, 11.495565, 11.510744, 11.573912, 11.692603, 11.867609, 12.097741, 12.376502, 12.69445, 13.03909, 13.396171, 13.75286, 14.132723, 14.456619, -999.0, 15.013323, 15.232368, 15.403331, 15.524743, 15.598823, 15.628752, 15.621209, 15.583071, 15.522541, 15.448029, 15.367778, 15.28981, 15.221546, 15.169065, 15.137166, 15.127272, 15.140369, 15.175196, 15.229729, 15.300282, 15.381946, 15.470299, 15.561097, 15.650753, 15.737549, 15.820256, 15.89977, 15.977968, 16.057486, 16.141966, 16.234447, 16.338512, 16.45688, 16.591022, 16.741774, 16.909342, 17.093513, 17.293243, 17.505873, 17.7295, 17.962448, 18.20347, 18.451479, 18.70529, 18.963926, 19.22663, 19.492228, 19.759706, 20.027353, 20.293968, 20.558214, 20.818615, 21.07407, 21.32338, 21.565083, 21.797686, 22.01867, 22.225426, 22.41473, 22.582762, 22.72577, 22.839725, 22.92058, 22.964596, 22.968102, 22.928932, 22.845785, 22.718346, 22.548262, 22.337759, 22.091785, 21.815985, 21.518143, 21.207327, 20.893145, 20.585968, 20.296608, 20.034988, 19.810814, 19.630877, 19.500755, 19.42375, 19.40029, 19.427896, 19.500042, 19.608143, 19.741219, 19.887594, 20.037558, 20.196207, 20.326075, 20.43564, 20.519577, 20.574635, 20.59912, 20.595442, 20.567307, 20.5194, 20.45711, 20.38583, 20.310804, 20.236683, 20.166815, 20.10367, 20.04784, 19.998869, 19.95572, 19.91672, 19.879734, 19.842653, 19.803627, 19.763025, 19.721916, 19.68286, 19.649632, 19.626081, 19.616644, 19.62592, 19.658407, 19.718561, 19.80962, 19.934124, 20.09371, 20.288366, 20.51758, 20.77817, 21.06681, 21.378939, 21.70953, 22.053518, 22.40552, 22.76002, 23.111301, 23.453466, 23.781301, 24.089788, 24.375544, 24.636316, 24.869823, 25.074242, 25.247845, 25.38947, 25.497707, 25.571743, 25.611732, 25.621292, 25.606754, 25.572126, 25.517796, 25.444826, 25.35761, 25.26157, 25.163347, 25.070078, 24.98725, 24.918278, 24.865683, 24.830368, 24.812283, 24.809757, 24.82014, 24.840048, 24.864958, 24.890722, 24.912823, 24.927113, 24.92982, 24.917315, 24.886148, 24.833086, 24.755146, 24.650501, 24.51708, 24.35369, 24.159388, 23.934849, 23.682276, 23.405104, 23.109516, 22.801977, 22.490448, 22.18288, 21.886822, 21.60935, 21.35688, 21.13505, 20.948664, 20.800472, 20.69338, 20.628456, 20.606455, 20.630045, 20.690819, 20.782911, 20.898039, 21.031044, 21.183357, 21.355082, 21.536083, 21.713194, 21.877981, 22.02549, 22.152706, 22.260654, 22.34966, 22.416925, 22.459616, 22.478796, -999.0, 22.459286, 22.42853, 22.3889, 22.342585, 22.291714, 22.238966, 22.187132, 22.138834, -999.0, 22.062841, 22.040018, 22.03067, 22.037926, 22.065071, 22.115015, 22.190336, 22.29175, 22.41723, 22.563353, 22.723465, 22.891222, 23.065517, 23.246775, 23.429888, 23.604856, 23.762012, 23.89206, 23.986021, 24.036503, 24.036308, 23.976835, 23.849478, 23.652582, -999.0, 23.2482, 22.923779, 22.573315, 22.209267, 21.838604, 21.468277, 21.106936, 20.763721, 20.448992, 20.173967, 19.948473, 19.779291, 19.671066, 19.620674, 19.623102, 19.671213, 19.756481, 19.8725, 20.01493, 20.177835, 20.352016, 20.52873, 20.70275, 20.869759, 21.023693, 21.157833, 21.26888, 21.359688, 21.432293, 21.485725, -999.0, 21.534863, 21.539936, 21.539562, 21.539322, 21.544819, 21.56168, 21.59552, 21.650427, 21.729914, 21.838251, 21.97915, 22.154552, 22.359743, 22.588802, 22.83373, 23.085968, 23.342108, 23.602497, 23.863998, 24.143883, 24.385136, 24.613113, 24.826767, 25.01908, 25.18089, 25.307894, 25.401308, 25.46184, -999.0, 25.498426, 25.483976, 25.45546, 25.418612, 25.379211, 25.343163, 25.31616, 25.303965, 25.310518, -999.0, 25.392443, 25.47083, 25.574461, 25.701057, 25.847986, 26.010265, 26.182455, 26.358809, 26.533392, 26.700521, 26.854671, 26.990395, 27.103563, -999.0, 27.248436, 27.276627, 27.275436, 27.247131, 27.194412, 27.121672, 27.033688, 26.936506, 26.836557, 26.740654, 26.655806, 26.588194, 26.542788, 26.524134, 26.53494, 26.577654, 26.652624, 26.759214, 26.894478, 27.05286, 27.227236, 27.408123, 27.587095, 27.760698, 27.926325, 28.080456, 28.219677, 28.341501, 28.44401, 28.52411, 28.57681, 28.59729, 28.586355, 28.547401, -999.0, 28.41641, -999.0, 28.261145, 28.17819, 28.093378, 28.008442, 27.927114, 27.854134, 27.792349, 27.742067, -999.0, 27.675932, 27.658258, 27.649008, 27.646448, 27.649143, 27.655933, 27.665628, -999.0, 27.690699, 27.705421, 27.721853, 27.740746, 27.76333, -999.0, 27.822708, 27.860712, 27.905884, 27.959518, 28.021288, 28.090027, 28.164972, 28.245499, 28.33987, 28.430037, 28.523144, 28.616547, 28.707592, 28.796179, 28.88321, 28.966341, 29.039011, 29.095224, 29.133942, 29.155212, 29.161581, 29.157158, 29.143633, 29.12026, 29.08693, 29.045252, 28.997255, 28.94675, 28.898218, 28.85449, 28.817049, -999.0, 28.768003, 28.759226, 28.761452, 28.774595, 28.798613, 28.833208, 28.877333, -999.0, 28.985193, 29.044895, 29.105848, 29.165497, 29.220978, 29.269426, 29.307978, -999.0, -999.0, 29.344118, 29.32974, 29.297705, 29.246143, 29.172054, 29.07312, 28.954395, 28.823927, 28.687996, 28.552227, 28.422485, 28.303493, 28.199415, 28.112028, 28.042637, 27.994661, 27.972563, 27.979158, -999.0, 28.076958, 28.16563, 28.277756, -999.0, -999.0, 28.7041, 28.85589, 29.002142, 29.136877, 29.254128, 29.349178, 29.417723, 29.456167, 29.462168, 29.434074, 29.3729, 29.280003, 29.1591, 29.014473, 28.850792, 28.673342, 28.48763, 28.299534, 28.114967, 27.939348, 27.7781, 27.63523, 27.51398, -999.0, 27.344078, 27.296589, 27.27328, 27.272964, 27.292807, 27.329344, 27.379412, 27.439829, 27.506962, 27.57702, 27.646461, 27.71369, 27.777899, 27.839685, 27.900085, 27.957043, 28.005232, 28.040668, 28.063932, 28.076313, 28.08122, 28.08279, 28.082094, 28.077446, 28.06585, 28.047888, 28.022106, 27.990095, 27.953503, 27.911385, 27.861866, -999.0, 27.737896, 27.662382, 27.576458, 27.479496, 27.37334, 27.260551, 27.141735, 27.015482, 26.87918, 26.729326, 26.562822, 26.384018, -999.0, 26.109026, 25.93554, -999.0, 25.63588, 25.494467, 25.357985, 25.236183, 25.134378, 25.053682, 24.996014, 24.964136, 24.96089, 24.988297, 25.047777, 25.139555, 25.261665, 25.413908, -999.0, 25.802757, 26.02697, 26.254799, 26.474627, 26.674633, 26.843779, 26.975084, 27.060621, 27.093016, 27.065922, 26.980717, 26.844053, 26.659275, 26.428606, 26.156202, 25.853958, 25.534843, -999.0, 24.897978, 24.606594, 24.349068, 24.135769, 23.972084, 23.86348, 23.814432, 23.828747, 23.906582, 24.04407, 24.235504, 24.469994, 24.736761, -999.0, 25.32724, 25.629375, 25.920523, 26.18949, 26.426264, 26.62096, 26.766998, 26.8586, 26.895454, 26.879625, 26.813772, 26.702631, 26.55155, 26.369148, 26.165148, 25.952574, 25.745049, 25.550955, 25.37495, 25.221312, 25.092, 24.98947, 24.916035, 24.873796, 24.861105, 24.874098, 24.907656, -999.0, 25.01092, 25.073538, 25.140352, -999.0, 25.242092, 25.294203, 25.334915, 25.36263, 25.37726, 25.379473, 25.370384, 25.351915, 25.326479, 25.296997, 25.265734, 25.232662, 25.197412, 25.161211, 25.126085, 25.093842, 25.06606, 25.044064, 25.027569, 25.016209, 25.009754, 25.007889, 25.01014, 25.015818, 25.024084, 25.033937, -999.0, 25.055075, 25.06553, 25.075228, 25.083632, 25.090551, 25.096348, 25.101154, 25.10468, 25.10674, 25.10839, 25.111212, 25.116316, 25.124542, 25.136925, 25.154776, 25.179367, 25.211105, 25.25007, -999.0, 25.34916, 25.408476, 25.473183, 25.54231, 25.61382, 25.685186, 25.752953, 25.813295, 25.864244, -999.0, 25.938797, 25.960918, 25.971428, 25.970743, 25.959766, 25.939247, 25.910385, 25.875357, 25.83787, 25.801256, 25.765982, 25.731808, 25.698751, 25.666767, 25.636341, 25.60869, 25.58478, 25.564386, 25.54707, 25.531937, 25.517765, 25.503653, 25.489017, 25.473173, 25.455797, -999.0, 25.42706, 25.407925, 25.390373, 25.375082, 25.362583, 25.3531, 25.346764, 25.344288, 25.346806, 25.354982, 25.370165, 25.389435, 25.413885, 25.443382, 25.476524, 25.511179, 25.545635, 25.57837, 25.607637, 25.631405, -999.0, 25.655247, 25.652962, 25.639652, 25.614458, 25.576681, 25.527628, 25.469372, 25.406794, 25.345362, 25.287195, 25.232328, 25.182274, 25.139688, 25.10661, 25.083162, -999.0, 25.068619, 25.082644, 25.111338, 25.14969, 25.192425, 25.234083, 25.269926, 25.30053, 25.327581, 25.347765, 25.355131, 25.347258, 25.32749, 25.298227, 25.259596, 25.211897, 25.157915, 25.101631, -999.0, 24.99364, 24.946129, 24.905043, 24.871698, -999.0, 24.838675, 24.830055, 24.834742, 24.854673, 24.886396, 24.923298, 24.960468, 24.994387, 25.021456, 25.039478, 25.046373, -999.0, 25.02002, 24.984554, 24.934113, 24.869217, 24.792366, 24.70634, 24.61358, 24.516186, 24.414621, 24.308634, 24.200008, 24.092924, -999.0, 23.89912, 23.814795, 23.732742, 23.643671, 23.544846, 23.440178, 23.33183, 23.21863, 23.099155, -999.0, 22.82632, 22.665585, 22.48749, 22.293282, 22.090076, 21.884544, -999.0, 21.578081, 21.379509, 21.190844, 21.016884, 20.860912, 20.726025, 20.614552, 20.52691, 20.462755, 20.418436, 20.3881, 20.372826, 20.36482, -999.0, 20.35683, -999.0, 20.335175, 20.309248, 20.269058, 20.211466, 20.13438, 20.036144, 19.91643, 19.77638, 19.617126, 19.440653, 19.249014, 19.044298, 18.828571, 18.604237, 18.373821, 18.139484, 17.902834, 17.665707, 17.429083, 17.193752, 16.958576, 16.721409, 16.481201, -999.0, 15.991999, 15.744115, -999.0, 15.242143, 14.984813, 14.724368, 14.463809, 14.203261, 13.940909, 13.676744, 13.416396, 13.165651, 12.926332, 12.698842, 12.483127, -999.0, 12.083427, 11.900729, 11.7313795, 11.575656, 11.433828, 11.306218, -999.0, 11.090835, 10.998472, -999.0, 10.837281, 10.773363, 10.722743, 10.686213, 10.664337, 10.656483, 10.661623, 10.67773, 10.702758, 10.736376, 10.77901, 10.830628, -999.0, 10.956962, 11.026584, 11.096172, 11.164088, 11.228817, 11.28798, 11.338931, 11.379495, 11.408205, 11.423873, 11.42631, -999.0, 11.390744, 11.350624, 11.294668, 11.223495, 11.137867, 11.040274, 10.932511, 10.8152485, 10.688915, 10.55596, -999.0, 10.353701, 10.224387, 10.106386, 10.003539, 9.9171505, 9.848443, 9.796455, 9.759987, 9.737466, 9.726985, 9.727243, 9.736402, 9.751947, 9.771261, 9.791429, 9.809405, 9.82224, 9.829138, -999.0, 9.826394, 9.819364, 9.8108, 9.802639, 9.796839, 9.795905, -999.0, 9.820466, 9.853117, 9.903029, 9.97051, 10.056055, 10.159373, 10.279929, 10.4161005, -999.0, 10.725578, 10.892752, 11.06372, 11.235518, 11.4051485, 11.570585, 11.730361, 11.884433, 12.03369, 12.177522, 12.313498, 12.439927, 12.557712, 12.667957, 12.77067, 12.865584, 12.95291, 13.033237, 13.107233, 13.175373, 13.237758, 13.293017, 13.339481, 13.377591, 13.40939, 13.43631, 13.459005, 13.47809, 13.4937315, 13.505967, 13.515075, 13.521451, 13.525599, 13.528328, 13.530575, -999.0, 13.538485, 13.546124, 13.557114, 13.571958, 13.590776, 13.613549, 13.639598, 13.668226, 13.699054, 13.731817, -999.0, 13.782632, 13.815101, 13.844007, 13.867174, 13.883809, 13.895092, 13.902217, 13.907606, 13.913746, 13.923891, 13.941636, 13.971118, 14.017175, 14.084682, 14.178402, 14.304549, 14.467427, 14.669858, 14.905771, 15.16467, 15.443534, 15.746352, 16.074219, 16.419888, 16.775806, 17.134905, 17.48943, 17.8331, 18.16184, 18.471199, 18.758726, 19.022472, 19.264122, -999.0, 19.691755, 19.87998, 20.051628, 20.206203, 20.34243, 20.458185, 20.55058, 20.623034, 20.66184, 20.678432, 20.678959, 20.665134, 20.632973, 20.58009, 20.512316, 20.437033, 20.361359, 20.293123, 20.23877, 20.201992, 20.186514, 20.19417, 20.226658, 20.286577, 20.376526, 20.495724, 20.639973, 20.806274, 20.993532, 21.199684, 21.416725, 21.634764, 21.846167, 22.044502, 22.223434, -999.0, 22.504364, 22.598017, 22.655622, 22.675404, 22.656658, 22.599646, -999.0, 22.38154, 22.228605, 22.053211, 21.86141, 21.659836, 21.455786, 21.25703, 21.07052, 20.901657, 20.755781, 20.63739, 20.550797, 20.498827, 20.483173, 20.504951, 20.56306, 20.656313, 20.780937, 20.932762, 21.106325, 21.295328, 21.493456, 21.694124, 21.890476, 22.076015, 22.244099, 22.390614, 22.512224, 22.607885, 22.679115, 22.727707, 22.75727, 22.771572, 22.774267, 22.769243, 22.75932, 22.74645, 22.731476, 22.713041, 22.690046, 22.660763, 22.62324, 22.575285, 22.514513, 22.439106, 22.348469, 22.24296, 22.126528, 22.003042, 21.877754, 21.756441, 21.645828, 21.553406, 21.486357, 21.450945, 21.453045, 21.494183, 21.575264, 21.69437, 21.847298, 22.027822, 22.22641, 22.433746, 22.64161, 22.84346, 23.036703, 23.236078, 23.393885, 23.51475, 23.594467, 23.643589, 23.670225, 23.67998, 23.678278, 23.668879, 23.653748, 23.63416, 23.610928, 23.58488, 23.557343, 23.530296, 23.504854, -999.0, 23.46198, 23.442097, 23.422277, 23.404879, 23.392925, 23.390425, 23.399961, 23.418505, 23.440264, 23.461357, 23.479996, 23.494463, 23.505016, 23.513535, 23.52574, 23.548714, -999.0, 23.644724, 23.72362, 23.825367, 23.950804, 24.099188, 24.268732, 24.452774, 24.641468, 24.822205, 24.979572, 25.100567, 25.180119, 25.214617, -999.0, 25.146969, -999.0, 24.906544, 24.727379, 24.513964, 24.271358, 24.01241, 23.752956, 23.511482, -999.0, 23.150938, 23.0456, 22.993343, -999.0, 23.050482, 23.16203, 23.330936, 23.553286, -999.0, 24.118689, 24.441952, 24.778833, 25.119982, -999.0, -999.0, 25.916756, 26.174427, 26.381994, 26.53465, 26.629599, 26.668087, 26.651655, 26.583683, 26.4684, -999.0, 26.22489, 26.029593, -999.0, 25.612814, 25.41459, 25.237751, 25.092161, -999.0, 24.92328, 24.904152, 24.933435, 25.00773, -999.0, 25.29288, 25.495466, 25.735722, 26.015066, 26.3277, 26.652788, 26.96877, 27.264454, -999.0, 27.768454, 27.971855, 28.138268, 28.259705, 28.33344, 28.372225, 28.39051, -999.0, 28.386923, 28.360434, 28.31656, -999.0, 28.189772, 28.11469, 28.03649, 27.956362, 27.876595, 27.802008, -999.0, 27.712568, 27.676159, -999.0, 27.681799, 27.733023, -999.0, 27.924818, 28.055237, 28.203592, 28.363613, -999.0, 28.598131, 28.732244, 28.835548, -999.0, -999.0, 28.891373, 28.817049, 28.69589, 28.528938, 28.317953, 28.066498, 27.782608, 27.473915, -999.0, 26.79865, 26.445946, -999.0, -999.0, 25.489616, -999.0, 25.060705, 24.936388, 24.882204, 24.904678, 25.00217, 25.161026, 25.365993, 25.60095, -999.0, 26.111929, 26.385082, -999.0, 26.953693, 27.233845, 27.492468, 27.71329, 27.884165, 27.994791, 28.04402, -999.0, -999.0, -999.0, 27.849333, 27.727818, 27.59338, 27.456078, 27.328926, 27.22427, 27.149746, 27.111172, 27.109997, -999.0, -999.0, 27.255463, 27.36592, 27.503868, 27.669388, 27.858479, 28.05914, 28.259594, -999.0, -999.0, -999.0, 28.886385, 29.034554, -999.0, 29.286234, -999.0, 29.497738, 29.598036, 29.68811, -999.0, 29.79283, -999.0, 29.862808, 29.884417, 29.888456, 29.870377, 29.822441, -999.0, 29.62143, -999.0, 29.292072, 29.09355, -999.0, 28.635015, 28.373596, -999.0, 27.818283, 27.532995, 27.244055, 26.953154, 26.663166, 26.386347, 26.144463, 25.949818, 25.790129, 25.651209, 25.527546, 25.416489, 25.318874, 25.239014, 25.178648, 25.135057, -999.0, 25.09746, 25.09332, 25.107874, -999.0, 25.195925, 25.27246, 25.373789, -999.0, 25.651678, 25.824736, 26.01441, -999.0, 26.420315, 26.62319, 26.81528, 26.987568, 27.135311, 27.258888, 27.35787, 27.429373, 27.470798, 27.484089, 27.473272, 27.447037, -999.0, 27.400953, 27.410715, 27.460957, -999.0, 27.73401, 27.966734, 28.25316, 28.583755, -999.0, -999.0, 29.752958, 30.17263, 30.600393, 31.037151, 31.465755, -999.0, 32.019287, 32.29035, 32.46271, 32.532257, -999.0, -999.0, 32.24514, 32.033466, -999.0, 31.513073, 31.224085, 30.927294, 30.632168, 30.350597, 30.09374, 29.868185, 29.678818, 29.526527, 29.409569, 29.325447, 29.266748, 29.241499, -999.0, 29.27234, 29.326868, 29.404083, 29.500784, 29.613316, 29.741251, 29.890072, 30.063244, 30.253307, 30.450472, -999.0, 30.857853, 31.065151, 31.263464, 31.444906, 31.609175, 31.756578, 31.881329, -999.0, 32.008965, 32.051624, 32.062534, 32.047543, 32.014545, 31.970419, 31.920782, 31.870897, 31.8255, 31.78911, 31.765076, 31.756218, 31.763536, -999.0, 31.823505, 31.872248, -999.0, 31.99197, 32.054783, 32.112972, 32.160824, 32.19421, 32.21134, 32.21027, 32.187794, 32.141174, 32.073654, 31.991398, 31.90042, 31.806541, 31.712244, -999.0, 31.501163, 31.379522, -999.0, 31.115055, 30.978401, 30.844501, 30.720297, 30.612038, -999.0, -999.0, -999.0, -999.0, -999.0, 30.35818, -999.0, 30.396889, 30.43934, -999.0, 30.562107, 30.636736, 30.716213, 30.797585, -999.0, -999.0, 31.033224, 31.101114, -999.0, -999.0, 31.239792, 31.26027, 31.26644, 31.259144, -999.0, 31.212559, 31.175943, -999.0, 31.08562, 31.040913, 30.99868, 30.956944, 30.914053, 30.868847, 30.820988, -999.0, 30.725716, 30.67729, 30.622225, 30.558681, 30.48815, 30.402973, -999.0, 30.219715, -999.0, 30.013763, 29.918152, -999.0, 29.785978, 29.759409, 29.762997, 29.799007, -999.0, 29.915737, -999.0, 30.167145, 30.326008, -999.0, 30.69444, 30.886505, 31.072489, 31.247112, 31.372513, 31.521952, -999.0, 31.783533, 31.88393, 31.957932, 32.005615, 32.02814, 32.030098, 32.01645, 31.990915, 31.956673, -999.0, 31.866528, 31.813017, 31.760263, 31.713308, 31.673752, 31.642496, 31.620573, 31.608727, -999.0, 31.617825, 31.640581, 31.67783, 31.731552, 31.801437, -999.0, 31.980902, 32.081776, -999.0, 32.295948, 32.415768, 32.54266, -999.0, 32.798447, 32.913864, 33.01194, -999.0, 33.14507, -999.0, -999.0, -999.0, -999.0, -999.0, 33.070526, 33.010185, 32.94511, 32.879196, -999.0, 32.760338, 32.715134, -999.0, 32.671886, 32.677265, 32.699303, -999.0, 32.796257, 32.872993, -999.0, 33.06674, 33.171272, -999.0, 33.315567, 33.398483, 33.46967, 33.529408, -999.0, 33.61931, 33.65007, 33.67202, -999.0, 33.69827, 33.70699, 33.71567, 33.726345, -999.0, -999.0, 33.788498, -999.0, 33.8721, 33.929317, 33.99508, 34.06606, 34.139713, 34.21412, 34.28713, 34.35652, 34.420193, 34.476917, 34.52591, -999.0, 34.59887, 34.624035, -999.0, 34.63671, 34.62175, 34.58778, 34.533394, 34.45831, -999.0, 34.24684, 34.114178, 33.970127, 33.81988, 33.66377, 33.500427, 33.32996, 33.15413, -999.0, -999.0, 32.659954, 32.5386, 32.453747, -999.0, 32.400005, -999.0, -999.0, -999.0, 32.65508, -999.0, -999.0, 33.13022, 33.302906, 33.468315, -999.0, -999.0, -999.0, 34.042862, 34.18027, 34.312214, 34.431183, 34.530266, 34.61278, 34.68539, 34.74741, 34.792656, -999.0, -999.0, 34.80749, 34.7752, -999.0, 34.663822, 34.589878, 34.508175, -999.0, -999.0, 34.30279, 34.237156, -999.0, -999.0, 34.15712, -999.0, 34.235985, 34.325687, -999.0, 34.511467, 34.661343, 34.824677, 34.999542, -999.0, 35.38342, 35.577103, -999.0, 35.933937, -999.0, -999.0, 36.336384, 36.460377, 36.549274, 36.595333, -999.0, 36.546524, 36.448814, 36.299755, -999.0, -999.0, -999.0, 35.44506, 35.153008, 34.858513, 34.564957, 34.27501, -999.0, 33.75439, -999.0, 33.39957, 33.291065, 33.23507, -999.0, -999.0, 33.25487, 33.330112, 33.429203, 33.54241, 33.6612, 33.779247, 33.90076, -999.0, -999.0, -999.0, 34.367695, -999.0, 34.580124, 34.657776, -999.0, 34.76208, 34.78796, -999.0, -999.0, 34.76183, -999.0, 34.630363, 34.528965, -999.0, 34.279716, 34.137646, -999.0, 33.80112, -999.0, -999.0, 33.297203, 33.107502, 32.947067, 32.81159, 32.697002, 32.60514, -999.0, -999.0, -999.0, -999.0, 32.50158, 32.54864, 32.61908, 32.705303, 32.800148, 32.898342, -999.0, 33.09495, 33.20008, 33.308548, 33.41233, 33.50583, 33.58669, 33.651794, -999.0, 33.728573, 33.738655, 33.730526, -999.0, 33.67137, -999.0, 33.617638, 33.59523, 33.592396, 33.61072, 33.652565, 33.721844, 33.823017, 33.9596, 34.133896, 34.343533, 34.578537, -999.0, 35.09865, -999.0, -999.0, 35.87792, -999.0, 36.24601, 36.366077, 36.43953, 36.46359, 36.43526, 36.352196, 36.216007, -999.0, 35.794353, 35.50622, 35.1635, 34.77543, -999.0, -999.0, 33.757366, 33.43291, 33.16963, 32.957108, 32.79562, 32.68661, 32.631065, 32.631516, 32.690823, -999.0, 32.886578, 33.077293, 33.292492, 33.51157, -999.0, -999.0, -999.0, 34.265305, 34.40894, 34.52482, 34.614403, -999.0, 34.685246, 34.684338, 34.66677, 34.639744, 34.611275, 34.587997, 34.57438, 34.574467, -999.0, 34.60038, 34.63112, 34.665558, 34.699825, 34.7382, 34.785095, 34.83602, -999.0, -999.0, -999.0, -999.0, 34.99612, -999.0, 35.037495, 35.058422, 35.08445, -999.0, 35.159332, 35.210545, 35.271732, -999.0, -999.0, 35.483192, 35.601727, 35.74706, 35.92047, 36.115944, 36.326023, 36.542126, 36.75716, 36.97673, 37.21194, -999.0, -999.0, -999.0, 38.081577, 38.297997, 38.484715, 38.639927, 38.760807, -999.0, -999.0, -999.0, -999.0, 38.893654, 38.8526, -999.0, 38.7217, 38.640327, 38.553776, 38.465763, -999.0, 38.307133, 38.250298, -999.0, 38.184013, 38.17045, 38.169823, 38.18148, 38.20349, 38.233936, 38.27198, 38.3172, 38.369972, 38.431164, -999.0, 38.5742, 38.651134, 38.73152, 38.816372, 38.905975, 39.000618, -999.0, -999.0, -999.0, 39.367188, 39.46927, 39.56464, 39.656647, 39.74674, 39.83089, -999.0, 39.968105, 40.021904, 40.069218, 40.099277, 40.115543, -999.0, 40.10521, 40.07837, 40.037064, -999.0, 39.914967, 39.841713, -999.0, 39.74065, -999.0, 39.662846, 39.65812, 39.672894, 39.70528, -999.0, 39.83655, -999.0, 40.049507, -999.0, 40.291115, 40.40266, -999.0, -999.0, -999.0, 40.72929, 40.77268, 40.801174, 40.81611, -999.0, 40.818993, 40.81277, 40.804802, -999.0, 40.798477, -999.0, 40.826538, 40.86164, -999.0, -999.0, 40.9956, 41.057842, 41.124733, 41.19842, -999.0, -999.0, 41.47062, -999.0, -999.0, 41.711056, -999.0, -999.0, 41.812454, 41.82352, -999.0, -999.0, 41.782673, 41.75327, 41.72068, 41.687473, 41.65607, 41.629246, -999.0, 41.61189, 41.63315, -999.0, -999.0, -999.0, 41.931694, -999.0, 42.173664, -999.0, 42.388184, 42.544987, -999.0, 42.84976, -999.0, 43.069992, 43.134613, 43.16835, -999.0, 43.150036, -999.0, -999.0, -999.0, 42.88004, 42.755615, 42.61998, 42.481625, -999.0, -999.0, -999.0, 42.046234, 41.97703, -999.0, 41.897865, -999.0, 41.901257, 41.93236, 41.98143, -999.0, 42.1196, 42.19999, -999.0, 42.329033, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 42.650753, 42.641655, -999.0, 42.604687, -999.0, -999.0, 42.484425, 42.43499, 42.38619, -999.0, 42.317802, -999.0, 42.29349, 42.297398, -999.0, -999.0, 42.369194, -999.0, 42.449005, 42.498062, -999.0, 42.607864, 42.662315, -999.0, 42.730244, 42.761177, -999.0, 42.77509, 42.753628, -999.0, -999.0, -999.0, 42.4989, -999.0, 42.29535, 42.176888, 42.06055, 41.98429, 41.991062, -999.0, -999.0, -999.0, 42.813484, -999.0, 42.9241, -999.0, 39.627464, -999.0, -999.0, -999.0, -999.0, -999.0, 4.802821, 1.2159203, 0.7654329, -999.0, -999.0, -999.0, -999.0, 0.93554544, 0.23260392, -999.0}
wdir =
  {197.0003, -999.0, -999.0, 195.6804, 195.74545, -999.0, -999.0, -999.0, 196.43236, 196.68898, 196.95229, 197.21811, 197.49294, 197.77861, 198.0711, 198.3688, 198.66895, 198.9682, 199.26196, 199.54472, 199.8133, 200.0666, 200.30177, 200.51367, 200.69691, 200.84904, 200.9682, 201.05284, 201.10252, 201.11609, 201.09395, 201.03813, 200.95735, 200.86209, 200.75932, 200.65384, 200.54836, 200.44218, 200.33601, 200.23494, 200.1446, 200.06877, 200.01033, 199.96814, 199.93718, 199.91504, 199.90259, 199.89973, 199.90126, 199.90074, 199.89372, 199.8772, 199.85075, 199.81807, 199.78174, 199.74068, 199.69362, 199.64165, 199.58652, 199.52959, 199.46829, 199.42151, 199.3992, 199.41644, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 202.37398, 203.0215, 203.75735, 204.5509, -999.0, 206.2177, -999.0, -999.0, -999.0, 209.86786, -999.0, 212.30573, -999.0, 215.46114, -999.0, 219.34543, 221.46535, 223.58272, -999.0, -999.0, -999.0, -999.0, -999.0, 230.05357, 229.49168, 228.5182, 227.2418, 225.77074, 224.20668, 222.6274, 221.08879, 219.62994, 218.27628, 217.04645, 215.95781, 215.02626, 214.26643, 213.67897, 213.2688, 213.03406, 212.97061, 213.07585, 213.3399, 213.7497, 214.27596, 214.88087, 215.51678, 216.12794, 216.66144, 217.07208, 217.31883, 217.37886, 217.24084, 216.92162, 216.4452, 215.84216, 215.14647, 214.38986, 213.60556, 212.81938, 212.05458, 211.32841, 210.65068, 210.0287, 209.47182, 208.99178, 208.60129, 208.31305, 208.13896, 208.0796, 208.13512, 208.31152, 208.61618, 209.05002, 209.60411, 210.26743, 211.02502, 211.8608, 212.76144, 213.71385, 214.69792, 215.68825, 216.66167, 217.60078, 218.49313, 219.34077, 220.22931, 221.00072, 221.73956, 222.44757, 223.12619, 223.77965, 224.41939, 225.05754, 225.70605, 226.3768, 227.07938, 227.82103, 228.60931, 229.45139, 230.35205, 231.30806, 232.3115, 233.3478, 234.39717, 235.44136, 236.46407, 237.44745, 238.36818, 239.20393, 239.93715, 240.5561, 241.06305, 241.47226, 241.78987, 242.00711, 242.11792, 242.13235, 242.06294, 241.91466, 241.689, 241.39024, 241.02655, 240.60371, 240.12227, 239.58212, 238.9902, -999.0, 237.6953, 237.01503, 236.32889, 235.65004, 234.99167, 234.36794, 233.79347, 233.283, 232.85152, 232.5141, 232.28261, 232.16911, 232.17969, 232.31897, 232.58926, 232.98991, 233.51953, 234.17194, 234.93695, 235.79103, 236.70642, 237.6557, 238.61038, 239.54305, 240.4292, 241.24399, 241.96483, 242.57204, 243.0582, 243.42047, 243.65556, 243.76187, 243.74197, 243.60551, 243.36064, 243.01273, 242.56702, 242.03726, 241.44308, 240.80705, 240.15472, 239.50514, 238.85619, 238.20515, 237.56866, 236.9707, 236.4289, 235.95605, 235.56348, 235.25662, 235.04147, 234.92668, 234.9204, 235.02155, -999.0, 235.52078, 235.91315, 236.39629, 236.95724, 237.58011, 238.2418, 238.91586, 239.64774, 240.28947, 240.8938, 241.44527, 241.9291, 242.33377, 242.64816, 242.86087, 242.96027, 242.93591, 242.78134, 242.49593, 242.09969, 241.61865, 241.08781, 240.54578, 240.0066, 239.4622, 238.91939, 238.41362, 237.98126, 237.64557, 237.42625, 237.33302, 237.3685, -999.0, 237.82657, -999.0, -999.0, 239.3898, 240.06883, 240.79337, 241.52707, 242.22395, 242.8587, 243.44182, 243.98376, 244.47812, 244.91531, 245.29199, 245.60855, 245.8658, 246.06494, 246.21086, 246.32104, 246.41408, 246.49875, -999.0, 246.66312, 246.76006, 246.87932, 247.0264, 247.2053, 247.41403, 247.64702, 247.8873, 248.10822, 248.2804, 248.37251, 248.35796, 248.22867, 247.98322, 247.62141, 247.14484, 246.56462, 245.90106, 245.17708, 244.42271, 243.66508, 242.92755, 242.22926, 241.58214, 240.9929, 240.4651, 239.99788, 239.58899, 239.22893, 238.90681, 238.60936, 238.3214, 238.02112, 237.6764, 237.25415, 236.72595, 236.06554, 235.25795, 234.29782, 233.19539, 231.97856, 230.68672, 229.37003, 228.08311, 226.8915, 225.85558, 225.01555, 224.51773, 224.07208, 223.84753, 223.84042, 224.04022, 224.43571, 225.01276, 225.83727, 226.74312, 227.77647, 228.91635, 230.12784, 231.37697, 232.63235, 233.8616, 235.02864, 236.09415, 237.02136, 237.7864, 238.36366, 238.7313, 238.86774, 238.75542, 238.38602, 237.7542, 236.87741, 235.77359, 234.4731, 233.01337, 231.44221, 229.81781, 228.2012, 226.65305, 225.23279, 223.98538, 222.95319, 222.16736, 221.64934, 221.40375, 221.41203, 221.65572, 222.10515, 222.73167, 223.50134, 224.37866, 225.32312, 226.29037, 227.24217, 228.14908, 228.98189, 229.71953, 230.34213, 230.8407, 231.21172, 231.45094, 231.55801, 231.53415, 231.39015, 231.13843, 230.79556, 230.38159, 229.91907, 229.43327, 228.951, 228.49835, 228.10252, 227.78714, 227.57434, 227.47987, 227.51572, 227.69807, 228.04593, 228.57431, 229.28394, 230.17438, 231.24364, 232.48547, 233.88118, 235.4049, 237.05396, 238.85492, 240.8152, 242.84555, 244.83548, 246.7328, 248.51967, 250.17685, 251.69864, 253.07732, 254.28925, 255.31082, 256.14044, 256.78668, 257.25662, 257.56604, 257.73178, 257.77927, -999.0, 257.61972, 257.439, 257.24442, 257.03546, 256.82968, 256.64307, 256.49033, 256.3735, 256.29193, 256.24756, 256.2434, 256.2878, 256.39697, 256.58395, 256.8532, 257.20804, 257.65436, 258.19864, 258.8487, 259.61282, 260.49506, 261.4836, 262.56778, 263.7257, 264.93304, -999.0, 267.36874, 268.5309, 269.61832, 270.6067, 271.47635, 272.2091, 272.79562, 273.22958, 273.50476, 273.6223, 273.58392, 273.41046, 273.12228, 272.74133, 272.28992, 271.77762, 271.20456, 270.57956, 269.92496, 269.26373, 268.6112, 267.98593, 267.4053, 266.88358, 266.4331, 266.0549, 265.75006, -999.0, 265.32214, 265.16953, 265.0317, 264.88824, 264.7198, 264.50912, 264.2476, 263.92288, 263.5246, 263.04233, 262.48123, 261.8598, 261.1943, 260.5093, 259.82965, 259.18405, 258.60422, 258.12515, 257.78598, 257.6274, 257.68552, 257.99863, 258.58173, 259.44965, 260.59314, 261.98907, 263.59952, 265.36548, 267.2234, 269.10236, 270.93182, 272.65717, 274.22894, 275.61563, 276.80106, 277.778, 278.56686, 279.18906, 279.69376, 280.13013, 280.54605, 280.99374, 281.53333, 282.22665, 283.12363, 284.24023, 285.59985, 287.23026, 289.1514, 291.3301, 293.68915, 296.15268, 298.63882, 301.06567, 303.35568, 305.4429, 307.28394, 308.85327, 310.1459, 311.26978, 312.03897, -999.0, 312.93607, 313.096, 313.07938, 312.899, 312.56854, 312.10178, 311.51596, 310.82602, 310.0433, 309.1793, 308.25165, 307.2816, 306.2982, 305.33875, 304.44083, 303.63736, 302.96164, 302.44257, 302.10587, 301.96783, 302.0365, 302.31537, 302.7979, 303.4759, 304.3311, 305.3447, 306.49335, 307.75, 309.07922, 310.4356, 311.776, 313.06055, 314.24887, 315.30136, 316.1803, 316.85583, 317.30548, 317.51428, 317.48138, 317.21027, 316.7196, 316.03152, 315.17645, 314.18845, 313.09894, 311.93854, 310.7384, 309.53384, 308.3586, 307.241, 306.20584, 305.2684, 304.43515, 303.71277, 303.10483, 302.61362, 302.2334, 301.95673, 301.7738, 301.67255, 301.6405, 301.66406, 301.73007, 301.82922, 301.95392, 302.10626, 302.29367, 302.524, 302.80753, 303.1555, 303.58118, 304.0997, 304.72968, 305.49167, 306.40378, 307.47974, 308.7275, 310.13956, 311.70416, 313.39954, 315.19724, 317.05737, 318.93222, 320.77438, 322.5379, 324.1813, 325.67172, 326.98166, 328.08997, 329.0562, 329.6957, 330.10748, 330.29495, 330.27005, 330.04178, 329.61765, 329.0054, 328.22333, 327.29544, 326.24435, 325.09366, 323.86816, 322.59238, 321.2914, 319.98572, 318.69394, 317.43146, 316.2092, 315.03455, 313.9063, 312.82214, 311.77887, 310.7734, 309.80588, 308.8786, 307.99188, 307.14438, 306.33633, 305.5738, 304.86444, 304.2202, 303.65512, 303.1795, 302.79947, 302.5194, 302.33664, 302.24646, 302.2365, 302.29257, 302.40204, 302.55203, 302.72705, 302.9081, 303.07852, 303.23096, 303.36017, 303.46613, 303.5525, 303.62216, 303.68143, 303.73862, 303.81345, 303.92984, 304.115, 304.39453, 304.76825, 305.21332, 305.7228, 306.3176, 307.0195, 307.8369, 308.77512, 309.81918, 310.935, 312.09225, 313.2612, 314.4095, 315.50665, 316.52216, 317.43103, 318.21313, 318.85388, 319.3507, 319.7011, 319.9135, 319.99768, 319.97388, 319.86673, 319.70233, 319.50977, 319.3178, 319.1519, 319.03796, 318.99405, 319.0373, 319.1803, 319.43094, 319.79437, 320.26508, 320.83606, 321.48776, 322.19614, 322.9306, 323.65506, 324.33487, 324.93857, 325.43552, 325.8053, 326.02747, 326.0906, 325.98856, 325.70023, 325.3082, 324.8292, 324.3052, 323.76416, 323.20715, 322.63968, 322.09735, 321.6205, 321.22888, 320.92813, 320.71786, 320.58505, 320.51883, 320.5158, 320.57352, 320.6838, -999.0, 321.0109, 321.18716, 321.34592, 321.48276, 321.59512, 321.68393, 321.75235, 321.80734, -999.0, 321.91525, 321.98184, 322.06415, 322.16864, 322.30237, 322.47464, 322.69513, 322.9651, 323.2751, 323.61365, 323.9647, 324.31332, 324.65225, 324.97644, 325.27615, 325.538, 325.7498, 325.90076, 325.9809, 325.98468, 325.9075, 325.7478, 325.50723, 325.19485, -999.0, 324.6436, 324.25995, 323.89844, 323.58304, 323.32062, 323.11914, 322.99323, 322.9587, 323.0231, 323.18668, 323.44055, 323.7621, 324.12933, 324.529, 324.94687, 325.3566, 325.7279, 326.0392, 326.27756, 326.43134, 326.49277, 326.45526, 326.31738, 326.08087, 325.75995, 325.3783, 324.95126, 324.48465, 323.98843, 323.48633, -999.0, 322.542, 322.10245, 321.69055, 321.3214, 321.00464, 320.73102, 320.49002, 320.2788, 320.09598, 319.93405, 319.78073, 319.6264, 319.46747, 319.30057, 319.12274, 318.93118, 318.72162, 318.4908, 318.24185, 317.9599, 317.70035, 317.42517, 317.12296, 316.80582, 316.49414, 316.1984, 315.92255, 315.6727, -999.0, 315.25955, 315.09003, 314.9351, 314.7939, 314.6688, 314.5564, 314.4453, 314.32587, 314.19458, -999.0, 313.88202, 313.6892, 313.46637, 313.21387, 312.93442, 312.6372, 312.33, 312.01263, 311.68356, 311.35098, 311.0299, 310.73032, 310.45535, -999.0, 309.99832, 309.8314, 309.71375, 309.65012, 309.6449, 309.7005, 309.81894, 309.9985, 310.23724, 310.53207, 310.87845, 311.26773, 311.687, 312.12463, 312.57117, 313.0166, 313.44757, 313.84967, 314.20865, 314.51062, 314.74408, 314.9037, 314.98636, 314.99826, 314.94775, 314.8431, 314.6921, 314.4978, 314.25806, 313.97388, 313.6545, 313.3084, 312.94022, 312.55533, -999.0, 311.80743, -999.0, 311.19122, 310.93253, 310.70483, 310.50815, 310.35104, 310.24594, 310.1944, 310.1843, -999.0, 310.26053, 310.3432, 310.44305, 310.54504, 310.63858, 310.7169, 310.77393, -999.0, 310.81342, 310.78973, 310.73245, 310.64172, 310.52185, -999.0, 310.2299, 310.0871, 309.96664, 309.88293, 309.842, 309.84503, 309.89514, 309.996, 310.16925, 310.3842, 310.65402, 310.97366, 311.33636, 311.7333, 312.1522, 312.5781, 312.99335, 313.38327, 313.7445, 314.07507, 314.37018, 314.62454, 314.83392, 314.9962, 315.11032, 315.17953, 315.20685, 315.19336, 315.14035, 315.0528, 314.9394, -999.0, 314.67255, 314.5399, 314.41788, 314.3115, 314.21854, 314.13205, 314.04932, -999.0, 313.9041, 313.84198, 313.78638, 313.74127, 313.7121, 313.70123, 313.70737, -999.0, -999.0, 313.76266, 313.78302, 313.80197, 313.81927, 313.83057, 313.83096, 313.81693, 313.78598, 313.74088, 313.68768, 313.62534, 313.54065, 313.4223, 313.27655, 313.11353, 312.9405, 312.7655, 312.59872, -999.0, 312.33228, 312.24542, 312.19336, -999.0, -999.0, 312.26523, 312.37094, 312.5184, 312.69888, 312.90323, 313.12463, 313.35715, 313.59802, 313.84775, 314.10632, 314.37106, 314.63736, 314.89343, 315.12622, 315.33133, 315.5092, 315.65784, 315.77475, 315.85797, 315.90695, 315.9205, 315.89603, 315.83102, -999.0, 315.5956, 315.4404, 315.26834, 315.08588, 314.90265, 314.7291, 314.57422, 314.44577, 314.34937, 314.28772, 314.26465, 314.2881, 314.3667, 314.50598, 314.70926, 314.9751, 315.29507, 315.66296, 316.07343, 316.52036, 316.99118, 317.47034, 317.94193, 318.39072, 318.84613, 319.2253, 319.56882, 319.86646, 320.10693, 320.28516, 320.39905, -999.0, 320.44403, 320.38895, 320.29233, 320.1633, 320.01743, 319.87228, 319.73935, 319.6263, 319.5472, 319.51926, 319.557, 319.65335, -999.0, 319.88165, 320.07504, -999.0, 320.53574, 320.81412, 321.11392, 321.40686, 321.67178, 321.8988, 322.07712, 322.20203, 322.27094, 322.28058, 322.2282, 322.1132, 321.93652, 321.69614, -999.0, 321.02795, 320.6221, 320.19858, 319.77774, 319.37708, 319.0061, 318.65793, 318.32684, 318.02048, 317.7497, 317.52496, 317.3574, 317.2514, 317.1968, 317.18506, 317.20724, 317.2528, -999.0, 317.36115, 317.3991, 317.4154, 317.40155, 317.34967, 317.25287, 317.10822, 316.91373, 316.66727, 316.36935, 316.02774, 315.66367, 315.29715, -999.0, 314.61795, 314.3276, 314.0782, 313.87555, 313.72574, 313.63593, 313.61224, 313.65933, 313.76825, 313.92593, 314.127, 314.37027, 314.6513, 314.95944, 315.28287, 315.60788, 315.9186, 316.20163, 316.4469, 316.64978, 316.81622, 316.95084, 317.05307, 317.1216, 317.15668, 317.16003, 317.14056, -999.0, 317.10208, 317.1112, 317.15527, -999.0, 317.30753, 317.45596, 317.64563, 317.87653, 318.14618, 318.45132, 318.7868, 319.14447, 319.51416, 319.8816, 320.23267, 320.55826, 320.8499, 321.1004, 321.3042, 321.45694, 321.5577, 321.60617, 321.60568, 321.5599, 321.4724, 321.34714, 321.1896, 321.00717, 320.80682, 320.59613, -999.0, 320.17368, 319.97867, 319.80838, 319.67377, 319.57938, 319.52036, 319.49442, 319.5052, 319.55652, 319.64584, 319.76727, 319.91214, 320.06924, 320.23288, 320.40738, 320.5949, 320.78232, 320.9529, -999.0, 321.21506, 321.30203, 321.36157, 321.39688, 321.41327, 321.4158, 321.40405, 321.3752, 321.33282, -999.0, 321.24637, 321.21478, 321.19516, 321.1856, 321.18298, 321.1921, 321.22302, 321.27896, 321.35135, 321.43246, 321.5226, 321.62375, 321.73694, 321.8632, 322.00055, 322.1423, 322.2827, 322.4189, 322.5484, 322.6675, 322.77203, 322.85605, 322.91257, 322.93707, 322.93182, -999.0, 322.8727, 322.80084, 322.7065, 322.59695, 322.47836, 322.3492, 322.20578, 322.05307, 321.904, 321.76953, 321.64474, 321.55563, 321.48328, 321.41986, 321.36465, 321.3193, 321.28015, 321.2396, 321.19293, 321.1434, -999.0, 321.04697, 320.99945, 320.9493, 320.89233, 320.82706, 320.7594, 320.69525, 320.6403, 320.60126, 320.58597, 320.6021, 320.65424, 320.74182, 320.86533, 321.02783, -999.0, 321.48453, 321.78375, 322.12482, 322.49304, 322.87918, 323.28278, 323.70157, 324.12192, 324.52808, 324.91495, 325.28387, 325.62952, 325.938, 326.1979, 326.4096, 326.57507, 326.69092, 326.752, -999.0, 326.69583, 326.5719, 326.38162, 326.12686, -999.0, 325.67242, 325.35977, 325.05203, 324.75604, 324.48077, 324.23404, 324.0225, 323.85126, 323.72513, 323.6447, 323.6106, -999.0, 323.66556, 323.74008, 323.83197, 323.93243, 324.03806, 324.14526, 324.25006, 324.3487, 324.43677, 324.50903, 324.55862, 324.58, -999.0, 324.5351, 324.4846, 324.41995, 324.341, 324.2519, 324.16138, 324.0779, 324.00677, 323.9536, -999.0, 323.89996, 323.8937, 323.89532, 323.902, 323.91147, 323.91953, -999.0, 323.90317, 323.85626, 323.7754, 323.65527, 323.49048, 323.27777, 323.02402, 322.7443, 322.4479, 322.13547, 321.77463, 321.43875, 321.10373, -999.0, 320.48752, -999.0, 320.02017, 319.85968, 319.75012, 319.69278, 319.6876, 319.7318, 319.81677, 319.93335, 320.08572, 320.2948, 320.57632, 320.91312, 321.2824, 321.6699, 322.06137, 322.44254, 322.80936, 323.16562, 323.5262, 323.90665, 324.28445, 324.6172, 324.86313, -999.0, 324.9931, 324.9198, -999.0, 324.64343, 324.38785, 324.04135, 323.61383, 323.1058, 322.51907, 321.86353, 321.17316, 320.4895, 319.8288, 319.19485, 318.58887, -999.0, 317.42633, 316.87112, 316.3417, 315.83798, 315.35977, 314.90732, -999.0, 314.05817, 313.63138, -999.0, 312.71487, 312.2466, 311.78183, 311.32544, 310.88422, 310.4668, 310.08264, 309.74094, 309.45078, 309.21414, 309.03015, 308.89386, -999.0, 308.72314, 308.67136, 308.63037, 308.58167, 308.50256, 308.36566, 308.14255, 307.81995, 307.40543, 306.89542, 306.27295, -999.0, 304.65555, 303.697, 302.66846, 301.59692, 300.5092, 299.43042, 298.38693, 297.399, 296.48602, 295.6728, -999.0, 294.70673, 294.28214, 294.07065, 294.0706, 294.24112, 294.54932, 294.97113, 295.47623, 296.02637, 296.58417, 297.18488, 297.71115, 298.20032, 298.6263, 298.96683, 299.21158, 299.35168, 299.3945, -999.0, 299.24966, 299.1044, 298.94147, 298.7815, 298.64597, 298.55228, -999.0, 298.54535, 298.64386, 298.8145, 299.05627, 299.36633, 299.73172, 300.13702, 300.5609, -999.0, 301.3754, 301.73236, 302.04016, 302.29633, 302.49747, 302.6373, 302.70966, 302.71692, 302.66864, 302.57834, 302.46613, 302.34802, 302.22473, 302.09537, 301.96158, 301.82462, 301.68414, 301.5385, 301.38596, 301.22595, 301.05865, 300.88943, 300.72546, 300.57327, 300.4396, 300.33118, 300.25244, 300.2068, 300.1904, 300.19766, 300.2216, 300.25385, 300.28635, 300.311, 300.31982, -999.0, 300.2495, 300.14365, 299.96835, 299.71274, 299.37424, 298.9565, 298.47693, 297.9486, 297.36798, 296.7304, -999.0, 295.7201, 295.0646, 294.44702, 293.87827, 293.36295, 292.89548, 292.47397, 292.10135, 291.78, 291.50815, 291.28342, 291.1045, 290.97, 290.87784, 290.82513, 290.80997, 290.83206, 290.8894, 290.9746, 291.07947, 291.20383, 291.35855, 291.55124, 291.7868, 292.07065, 292.40814, 292.80487, 293.2664, 293.79575, 294.39062, 295.04297, 295.75464, 296.54416, -999.0, 298.39008, 299.38766, 300.39514, 301.39456, 302.36588, 303.29233, 304.15906, 305.0385, 305.77182, 306.44095, 307.0424, 307.56808, 308.00168, 308.3271, 308.53278, 308.60675, 308.54108, 308.33087, 307.9714, 307.4639, 306.8173, 306.0582, 305.2116, 304.28363, 303.27817, 302.22324, 301.1606, 300.11185, 299.07104, 298.03836, 297.04352, 296.1183, 295.27667, 294.52393, 293.8641, -999.0, 292.8142, 292.41788, 292.10376, 291.87518, 291.73895, 291.6992, -999.0, 291.9019, 292.12946, 292.42682, 292.7875, 293.20477, 293.6644, 294.14542, 294.6262, 295.08588, 295.50317, 295.86533, 296.16092, 296.38058, 296.51843, 296.57184, 296.54663, 296.45056, 296.30084, 296.11636, 295.91602, 295.71875, 295.5397, 295.38882, 295.27536, 295.2032, 295.1759, 295.19296, 295.25223, 295.3487, 295.4748, 295.6246, 295.79468, 295.98163, 296.18353, 296.39798, 296.621, 296.8492, 297.08514, 297.3386, 297.61658, 297.92117, 298.2547, 298.6237, 299.03647, 299.50342, 300.0366, 300.6458, 301.33212, 302.09723, 302.93878, 303.8522, 304.8267, 305.8458, 306.8932, 307.9501, 308.9946, 309.99905, 310.9355, 311.78055, 312.51422, 313.12085, 313.58972, 313.90833, 314.0639, 314.04263, 313.84686, 313.43967, 312.916, 312.27435, 311.5299, 310.6911, 309.77103, 308.8012, 307.8159, 306.85162, 305.94815, 305.1406, 304.45834, 303.93274, 303.5863, 303.44168, 303.49942, -999.0, 304.17374, 304.73187, 305.40436, 306.18173, 307.04718, 307.95737, 308.8644, 309.721, 310.4803, 311.10605, 311.57385, 311.8593, 311.9462, 311.82224, 311.49698, 310.98737, -999.0, 309.51614, 308.61588, 307.64685, 306.6368, 305.6045, 304.56668, 303.54407, 302.5582, 301.6325, 300.789, 300.0361, 299.35275, 298.71634, -999.0, 297.5203, -999.0, 296.33932, 295.74103, 295.15414, 294.58987, 294.03903, 293.49246, 292.96616, -999.0, 292.08145, 291.75095, 291.50595, -999.0, 291.3005, 291.35596, 291.5283, 291.81293, -999.0, 292.65707, 293.19363, 293.7905, 294.4173, -999.0, -999.0, 295.93237, 296.473, 296.94284, 297.31317, 297.56342, 297.68173, 297.66138, 297.51492, 297.25464, -999.0, 296.68283, 296.2045, -999.0, 295.1223, 294.59195, 294.13577, 293.79385, -999.0, 293.5468, 293.65726, 293.95294, 294.3676, -999.0, 295.53387, 296.22598, 296.95422, 297.69153, 298.39478, 298.99222, 299.42203, 299.67197, -999.0, 299.6391, 299.3662, 298.92853, 298.32697, 297.5599, 296.63336, 295.5647, -999.0, 293.88, 292.84778, 291.94846, -999.0, 290.6368, 290.20258, 289.9083, 289.77414, 289.81714, 290.04163, -999.0, 290.69785, 291.27808, -999.0, 292.59695, 293.3159, -999.0, 294.7541, 295.41415, 296.0074, 296.51376, -999.0, 297.05887, 297.26035, 297.34183, -999.0, -999.0, 296.91254, 296.55557, 296.11557, 295.6136, 295.07477, 294.52197, 293.97205, 293.44022, -999.0, 292.4519, 292.012, -999.0, -999.0, 291.11902, -999.0, 290.98904, 291.0903, 291.3108, 291.65155, 292.0922, 292.58612, 293.09232, 293.5898, -999.0, 294.50925, 294.92865, -999.0, 295.70587, 296.06458, 296.37744, 296.62198, 296.79156, 296.88312, 296.8955, -999.0, -999.0, -999.0, 296.35632, 296.05283, 295.6905, 295.28296, 294.86383, 294.46674, 294.10608, 293.79004, 293.5222, -999.0, -999.0, 293.07562, 293.01578, 293.03403, 293.12344, 293.27722, 293.4867, 293.7413, -999.0, -999.0, -999.0, 294.69583, 294.9022, -999.0, 295.12265, -999.0, 295.01855, 294.8225, 294.51633, -999.0, 293.8591, -999.0, 293.0338, 292.51837, 292.03436, 291.594, 291.19608, -999.0, 290.5463, -999.0, 290.16324, 290.09302, -999.0, 290.1963, 290.35837, -999.0, 290.87714, 291.22214, 291.6157, 292.04926, 292.51184, 292.983, 293.43146, 293.83554, 294.20578, 294.55655, 294.89017, 295.205, 295.4996, 295.77167, 296.02118, 296.25223, -999.0, 296.56622, 296.7427, 296.8875, -999.0, 297.1138, 297.20554, 297.2835, -999.0, 297.37698, 297.382, 297.36298, -999.0, 297.25345, 297.14905, 297.01764, 296.87497, 296.72812, 296.57532, 296.4181, 296.26785, 296.1377, 296.04254, 295.99762, 296.00842, -999.0, 296.18637, 296.36, 296.57794, -999.0, 297.16003, 297.49573, 297.81726, 298.10086, -999.0, -999.0, 298.65247, 298.73303, 298.77148, 298.77838, 298.75607, -999.0, 298.65753, 298.54898, 298.41248, 298.24954, -999.0, -999.0, 297.59943, 297.35806, -999.0, 296.85562, 296.58853, 296.3146, 296.03732, 295.75867, 295.48206, 295.21622, 294.97192, 294.7605, 294.5935, 294.47864, 294.41464, 294.41452, -999.0, 294.58423, 294.75024, 294.96286, 295.20795, 295.46524, 295.72296, 295.98364, 296.24594, 296.4879, 296.68472, -999.0, 296.92053, 296.96146, 296.94983, 296.88257, 296.7524, 296.5544, 296.30597, -999.0, 295.8921, 295.60443, 295.3113, 295.01837, 294.7328, 294.46484, 294.22824, 294.03415, 293.88538, 293.78333, 293.7284, 293.72034, 293.75693, -999.0, 293.9474, 294.09326, -999.0, 294.45908, 294.65997, 294.8614, 295.05652, 295.2427, 295.4232, 295.5985, 295.75983, 295.8974, 296.01074, 296.10352, 296.1779, 296.23453, 296.27405, -999.0, 296.3059, 296.3008, -999.0, 296.25916, 296.2328, 296.21072, 296.1988, 296.20175, -999.0, -999.0, -999.0, -999.0, -999.0, 296.4987, -999.0, 296.7339, 296.87314, -999.0, 297.17966, 297.3421, 297.50647, 297.66913, -999.0, -999.0, 298.09836, 298.215, -999.0, -999.0, 298.4619, 298.49838, 298.51697, 298.52142, -999.0, 298.49628, 298.46252, -999.0, 298.3449, 298.2744, 298.2007, 298.1223, 298.03992, 297.95712, 297.87808, -999.0, 297.75, 297.6984, 297.6421, 297.5787, 297.5146, 297.45004, -999.0, 297.36176, -999.0, 297.30927, 297.2961, -999.0, 297.32004, 297.36218, 297.42645, 297.51584, -999.0, 297.70038, -999.0, 298.0137, 298.18402, -999.0, 298.51697, 298.66568, 298.79715, 298.9122, 298.9912, 299.07623, -999.0, 299.187, 299.20956, 299.2068, 299.17532, 299.11493, 299.03378, 298.94077, 298.84204, 298.74228, -999.0, 298.5304, 298.41397, 298.30453, 298.21603, 298.15744, 298.13596, 298.148, 298.18225, -999.0, 298.29306, 298.36288, 298.43546, 298.50598, 298.57428, -999.0, 298.70422, 298.75458, -999.0, 298.79266, 298.77502, 298.74042, -999.0, 298.66068, 298.626, 298.5957, -999.0, 298.5118, -999.0, -999.0, -999.0, -999.0, -999.0, 298.03702, 297.93707, 297.83997, 297.74323, -999.0, 297.55124, 297.46033, -999.0, 297.305, 297.2434, 297.19064, -999.0, 297.1257, 297.12302, -999.0, 297.1584, 297.18472, -999.0, 297.22064, 297.2411, 297.2595, 297.27225, -999.0, 297.26416, 297.2422, 297.2103, -999.0, 297.13226, 297.0896, 297.04343, 296.99377, -999.0, -999.0, 296.83954, -999.0, 296.7605, 296.7274, 296.70496, 296.70386, 296.72757, 296.77097, 296.82996, 296.90204, 296.9847, 297.07513, 297.17007, -999.0, 297.34738, 297.4205, -999.0, 297.48755, 297.47803, 297.43134, 297.34833, 297.23343, -999.0, 296.91214, 296.7068, 296.47772, 296.23187, 295.97678, 295.71854, 295.45047, 295.15674, -999.0, -999.0, 294.16785, 293.846, 293.53656, -999.0, 293.11584, -999.0, -999.0, -999.0, 292.3991, -999.0, -999.0, 292.2789, 292.33282, 292.423, -999.0, -999.0, -999.0, 293.09222, 293.37253, 293.69635, 294.03412, 294.35675, 294.66003, 294.94778, 295.21844, 295.4697, -999.0, -999.0, 296.14532, 296.36594, -999.0, 296.82385, 297.07272, 297.34415, -999.0, -999.0, 298.14584, 298.51117, -999.0, -999.0, 299.60034, -999.0, 300.21848, 300.4959, -999.0, 300.86005, 301.04282, 301.14774, 301.16992, -999.0, 301.02216, 300.88165, -999.0, 300.51462, -999.0, -999.0, 299.90735, 299.6772, 299.47226, 299.29474, -999.0, 299.05435, 299.00592, 299.00302, -999.0, -999.0, -999.0, 299.2556, 299.35468, 299.44168, 299.5145, 299.57428, -999.0, 299.64398, -999.0, 299.63797, 299.60165, 299.53842, -999.0, -999.0, 299.15256, 298.99554, 298.85272, 298.74014, 298.66833, 298.64786, 298.6801, -999.0, -999.0, -999.0, 299.16382, -999.0, 299.6546, 299.9487, -999.0, 300.59488, 300.92303, -999.0, -999.0, 301.66013, -999.0, 302.10446, 302.2595, -999.0, 302.40103, 302.3726, -999.0, 302.08444, -999.0, -999.0, 301.29138, 300.89288, 300.48117, 300.04608, 299.57715, 299.08493, -999.0, -999.0, -999.0, -999.0, 297.07755, 296.7877, 296.57877, 296.4409, 296.36877, 296.36337, -999.0, 296.55856, 296.758, 297.00858, 297.28143, 297.55713, 297.82806, 298.08444, -999.0, 298.49884, 298.6313, 298.70013, -999.0, 298.6325, -999.0, 298.43256, 298.25677, 298.0642, 297.8653, 297.67316, 297.5028, 297.36884, 297.277, 297.22778, 297.22217, 297.25797, -999.0, 297.44077, -999.0, -999.0, 297.87256, -999.0, 298.1686, 298.3158, 298.45508, 298.58096, 298.69138, 298.7845, 298.8566, -999.0, 298.91916, 298.89944, 298.83896, 298.73724, -999.0, -999.0, 298.33893, 298.1541, 297.94904, 297.70807, 297.4278, 297.11163, 296.77307, 296.43994, 296.1322, -999.0, 295.7178, 295.47922, 295.28735, 295.15268, -999.0, -999.0, -999.0, 294.99786, 294.9943, 294.9827, 294.95172, -999.0, 294.83005, 294.71674, 294.55145, 294.34848, 294.1347, 293.91287, 293.66016, 293.36572, -999.0, 292.8908, 292.57504, 292.259, 291.942, 291.63086, 291.3335, 291.05502, -999.0, -999.0, -999.0, -999.0, 290.06995, -999.0, 289.7493, 289.60184, 289.45602, -999.0, 289.1914, 289.07864, 288.97604, -999.0, -999.0, 288.74353, 288.6435, 288.52448, 288.37863, 288.2044, 288.00397, 287.7896, 287.57236, 287.34622, 287.09927, -999.0, -999.0, -999.0, 286.19678, 285.99298, 285.83746, 285.73834, 285.70407, -999.0, -999.0, -999.0, -999.0, 286.2921, 286.5549, -999.0, 287.16617, 287.4909, 287.81003, 288.11124, -999.0, 288.6189, 288.81393, -999.0, 289.06763, 289.11926, 289.11502, 289.05472, 288.94824, 288.80527, 288.63077, 288.42844, 288.2022, 287.9573, -999.0, 287.46222, 287.24835, 287.0696, 286.93207, 286.84213, 286.80463, -999.0, -999.0, -999.0, 287.0666, 287.21948, 287.39362, 287.59177, 287.81128, 288.0337, -999.0, 288.4267, 288.592, 288.74112, 288.83548, 288.8856, -999.0, 288.87515, 288.82114, 288.73456, -999.0, 288.4407, 288.23254, -999.0, 287.89227, -999.0, 287.44965, 287.24796, 287.06757, 286.91354, -999.0, 286.68408, -999.0, 286.54227, -999.0, 286.4652, 286.4499, -999.0, -999.0, -999.0, 286.49258, 286.49194, 286.47238, 286.43283, -999.0, 286.35535, 286.30023, 286.2418, -999.0, 286.1066, -999.0, 285.92743, 285.8235, -999.0, -999.0, 285.57605, 285.50085, 285.44196, 285.39792, -999.0, -999.0, 285.30698, -999.0, -999.0, 285.2202, -999.0, -999.0, 285.10336, 285.0338, -999.0, -999.0, 284.74118, 284.6184, 284.48828, 284.3537, 284.21216, 284.06012, -999.0, 283.7341, 283.57144, -999.0, -999.0, -999.0, 283.05365, -999.0, 282.90424, -999.0, 282.82736, 282.78598, -999.0, 282.72565, -999.0, 282.69843, 282.69373, 282.6933, -999.0, 282.70453, -999.0, -999.0, -999.0, 282.7875, 282.82233, 282.85544, 282.8825, -999.0, -999.0, -999.0, 282.90656, 282.90466, -999.0, 282.90494, -999.0, 282.9068, 282.90192, 282.88834, -999.0, 282.83704, 282.8017, -999.0, 282.73364, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 282.1417, 282.00122, -999.0, 281.80994, -999.0, -999.0, 281.56802, 281.5096, 281.4567, -999.0, 281.3961, -999.0, 281.3849, 281.39334, -999.0, -999.0, 281.50177, -999.0, 281.65903, 281.7543, -999.0, 281.96518, 282.07733, -999.0, 282.2487, 282.35675, -999.0, 282.53677, 282.613, -999.0, -999.0, -999.0, 282.87576, -999.0, 282.96564, 283.0009, 283.0318, 283.0591, 283.08215, -999.0, -999.0, -999.0, 283.13196, -999.0, 283.17004, -999.0, 283.19836, -999.0, -999.0, -999.0, -999.0, -999.0, 283.22876, 283.2406, 103.205414, -999.0, -999.0, -999.0, -999.0, 103.22321, 103.22102, -999.0}
dz =
  {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 3.6814237, 3.7369893, 3.8006434, 3.8703165, 3.9438467, 4.021242, 4.102512, 4.1854258, 4.267601, 4.3490386, 4.429741, 4.507741, 4.580894, 4.649195, 4.71264, 4.7699046, 4.819516, 4.8614645, 4.8957415, 4.921784, 4.9389524, 4.9472322, 4.9466085, 4.937248, 4.9193444, 4.892879, 4.8578334, 4.8149867, 4.765266, 4.708656, 4.645142, 4.5759315, 4.50249, 4.424813, 4.3428917, 4.2580705, 4.1720104, 4.084717, 3.9961905, 3.9075453, 3.820184, 3.7341177, 3.6493533, 3.5665205, 3.4864252, 3.4090774, 3.3344834, 3.2626693, 3.1936688, 3.1274908, 3.064137, 3.003046, 2.9434214, 2.885271, 2.8230147, 2.7668488, 2.7099922, 2.652444, 2.5942016, 2.5341668, 2.4712968, 2.4055867, 2.3370326, 2.2649047, 2.1885908, 2.1080806, 2.023364, 1.9345969, 1.8419294, 1.745348, 1.6448407, 1.5419238, 1.4381357, 1.3334767, 1.2279476, 1.1244675, 1.0260881, 0.93281955, 0.8446709, 0.7653171, 0.6986329, 0.64462954, 0.6033158, 0.57787114, 0.5717211, 0.58487195, -999.0, -999.0, -999.0, -999.0, -999.0, 1.0910197, 1.2463332, 1.4207178, 1.6141891, 1.8227422, 2.0417824, 2.27133, 2.5114174, 2.7568612, 3.0015955, 3.2456307, 3.4889877, 3.7268987, 3.9536493, 4.1692257, 4.3736205, 4.563612, 4.735274, 4.888556, 5.023429, 5.1386976, 5.232846, 5.3058243, 5.357588, 5.3888497, 5.4005327, 5.392604, 5.3650274, 5.3199196, 5.260042, 5.185387, 5.0959373, 4.9945173, 4.8848705, 4.767006, 4.6409144, 4.5095406, 4.3768597, 4.242896, 4.107653, 3.9736664, 3.8444211, 3.7199476, 3.6002545, 3.4870403, 3.382684, 3.287214, 3.2006412, 3.1235468, 3.056758, 3.000295, 2.954171, 2.917799, 2.8903167, 2.871728, 2.862043, 2.859895, 2.8632467, 2.8720844, 2.8864138, 2.9048305, 2.9252017, 2.9498415, 2.9742703, 2.9996724, 3.025023, 3.0503182, 3.0755541, 3.1008005, 3.126135, 3.1515574, 3.1770673, 3.2033808, 3.231297, 3.2608187, 3.2919486, 3.3253775, 3.361892, 3.4014976, 3.444199, 3.4901955, 3.5397165, 3.5927675, 3.649353, 3.7089732, 3.7710345, 3.8355396, 3.9024925, 3.9706573, 4.03854, 4.1061397, 4.1734595, 4.238734, 4.2997837, 4.3566017, 4.409187, 4.4558477, 4.494455, 4.524987, 4.547432, 4.560959, 4.5645065, 4.5580544, 4.5415854, 4.5155234, 4.480427, 4.4362826, 4.3830757, 4.3222747, 4.255847, 4.183797, 4.1061163, 4.0247965, 3.94255, 3.859391, 3.7753186, 3.6921804, 3.612545, 3.5364358, 3.46386, 3.3958821, 3.3340104, 3.2782671, 3.2286637, 3.1851861, 3.1478088, 3.1165414, 3.0913937, 3.0714867, 3.0555198, 3.0434854, 3.0353873, 3.029978, 3.025382, 3.0215793, 3.018568, 3.0152395, 3.009896, 3.0025136, 2.9930866, 2.9810345, 2.9654574, 2.9463377, 2.9236686, 2.8975704, 2.8682382, 2.8356702, 2.7998617, 2.7615087, 2.7217433, 2.680581, 2.6380222, 2.5949168, 2.5526707, 2.5113082, 2.4708333, 2.431767, 2.3949833, 2.360501, 2.328325, 2.2983556, 2.2704196, 2.2445173, 2.2206528, 2.1981466, 2.175809, 2.1514091, 2.1293857, 2.1063285, 2.080762, 2.052679, 2.022077, 1.9879905, 1.9491911, 1.9056685, 1.8574171, 1.8041464, 1.7454822, 1.6814182, 1.6119498, 1.5375253, 1.4587394, 1.3755937, 1.2880871, 1.197226, 1.1043617, 1.0095034, 0.9126553, 0.81508076, 0.71851814, 0.622982, 0.5284765, 0.43594894, 0.34672558, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 2.3769405, 2.5262573, 2.67893, 2.8346353, 2.9927397, 3.1532278, 3.3161075, 3.4972894, 3.6626287, 3.8285458, 3.9950495, 4.160771, 4.323732, 4.483925, 4.6413608, 4.794342, 4.9403634, 5.0794034, 5.2114615, 5.3349705, 5.4475594, 5.5491924, 5.639858, 5.7185497, 5.783742, 5.835382, 5.8734636, 5.897871, 5.908432, 5.9051113, 5.8878517, 5.8574963, 5.8153825, 5.7614946, 5.6958, 5.6198616, 5.536237, 5.4449434, 5.3459654, 5.2411666, 5.1336446, 5.02345, 4.9105873, 4.796731, 4.6846976, 4.5745482, 4.466296, 4.3611116, 4.26099, 4.165983, 4.0761085, 3.9919245, 3.9143925, 3.843541, 3.7793806, 3.7219393, 3.6712563, 3.6273396, 3.590197, 3.5595562, 3.534913, 3.51626, 3.5035996, 3.4966357, 3.4948163, 3.4981303, 3.5065782, 3.5200794, 3.5384822, 3.5617847, 3.5899885, 3.6232994, 3.6621127, 3.7064428, 3.756293, 3.81196, 3.8740187, 3.942492, 4.017387, 4.098777, 4.186801, 4.2814717, 4.3827987, 4.49041, 4.6035447, 4.722192, 4.846364, 4.9752073, 5.106949, 5.2415457, 5.3790092, 5.5181823, 5.656617, 5.794244, 5.9310713, 6.0659394, 6.1963563, 6.3222456, 6.443615, 6.5708065, 6.6787915, 6.7794385, 6.8727474, 6.9581156, 7.034588, 7.102132, 7.160724, 7.2103696, 7.251086, 7.282841, 7.3056006, 7.319999, 7.3271003, 7.326892, 7.319347, 7.3055425, 7.2873, 7.264634, 7.237532, 7.2071266, 7.175356, 7.1422515, 7.1078124, 7.072849, 7.0387664, 7.0055966, 6.9733477, 6.9423504, 6.913179, 6.8858476, 6.86036, 6.8367047, 6.814853, 6.794803, 6.776559, 6.7599735, 6.7447667, 6.7309384, 6.718491, 6.7072377, 6.6968293, 6.68726, 6.6785326, 6.67049, 6.662834, 6.6555614, 6.648673, 6.6421275, 6.635841, 6.6298127, 6.624045, 6.618686, 6.6140304, 6.610085, 6.606851, 6.6046677, 6.6042156, 6.605516, 6.60857, 6.613737, 6.6217527, 6.632645, 6.6464224, 6.6631756, 6.6830897, 6.706183, 6.732468, 6.76155, 6.792577, 6.825534, 6.860435, 6.896426, 6.9316382, 6.9660115, 6.9995484, 7.031251, 7.058911, 7.0824428, 7.101841, 7.1164217, 7.1246586, 7.126475, 7.121851, 7.1107836, 7.093291, 7.069351, 7.0389404, 7.0027447, 6.9624815, 6.918203, 6.869851, 6.818464, 6.7666545, 6.714527, 6.6620784, 6.6101465, 6.5607653, 6.513973, 6.469806, 6.428423, 6.3901505, 6.354992, 6.3229613, 6.2934613, 6.264972, 6.2374206, 6.2108235, 6.1841903, 6.1550593, 6.1232986, 6.088903, 6.0470414, 6.003333, 5.9541364, 5.8994355, 5.8389993, 5.7724056, 5.699625, 5.62064, 5.536219, 5.447858, 5.355584, 5.259391, -999.0, -999.0, -999.0, 4.848382, 4.740878, 4.6329556, 4.5246587, 4.415998, 4.307682, 4.201131, 4.096396, 3.9934871, 3.8926997, 3.7946317, 3.6993096, 3.6067412, 3.5171607, 3.431051, 3.3484325, 3.2693095, 3.1939924, 3.1231384, 3.0567734, 2.9949014, 2.9379292, 2.8867393, 2.8413665, 2.8018155, 2.768431, 2.7419736, 2.7224777, 2.7099495, 2.7044628, 2.7061768, 2.7151008, 2.7312489, 2.7543142, 2.7835798, 2.8190172, 2.8606386, 2.9078226, 2.9591, 3.0144145, 3.0737717, 3.1364715, 3.2008288, 3.2667696, 3.3342936, 3.4028127, 3.470899, 3.5384872, 3.605576, 3.6716418, 3.7353923, 3.796767, 3.855765, 3.9118319, 3.9635634, 4.0108886, 4.0538054, 4.091849, 4.123827, 4.149668, 4.169359, 4.1827884, 4.1896815, 4.1900115, 4.183763, 4.1712766, 4.1534753, 4.130404, 4.102056, 4.0690813, 4.033255, 3.9946778, 3.9533496, 3.9100301, 3.8668213, 3.8238473, 3.7811098, 3.7352695, 3.6966236, 3.6609654, 3.6282992, 3.599273, 3.5752118, 3.5561616, 3.5421305, 3.5332663, 3.529872, 3.5319667, 3.5395603, 3.552252, 3.5691774, 3.5903149, 3.6156714, 3.6445506, 3.675436, 3.7082753, 3.7430687, 3.7791986, 3.8153052, 3.8513339, 3.8872786, 3.9228616, 3.9574723, 3.991088, 4.023708, 4.055413, 4.086389, 4.1166472, 4.146191, 4.175262, 4.2044168, 4.233679, 4.263049, 4.2927365, 4.32323, 4.354545, 4.386678, 4.4196944, 4.4537635, 4.488894, 4.525089, 4.5622206, 4.599979, 4.638353, 4.6773467, 4.716731, 4.7559237, 4.7948995, 4.83366, 4.872096, 4.909925, 4.947133, 4.98372, 5.01972, 5.0552278, 5.0902534, 5.1248035, 5.1588354, 5.1922255, 5.2249746, 5.2570925, 5.2883124, 5.3178983, 5.3458104, 5.37205, 5.3962092, 5.4171615, 5.4348216, 5.449167, 5.4598465, 5.465923, 5.4673185, 5.464011, 5.455882, 5.442644, 5.4242735, 5.400764, 5.372239, 5.339069, 5.3012743, 5.2588525, 5.212056, 5.1616344, 5.1076255, 5.0500183, 4.9890623, 4.9255276, 4.8594575, 4.7908425, 4.7198086, 4.6467648, 4.5717406, 4.4947386, 4.41573, 4.334623, 4.2514105, 4.1660924, 4.078576, 3.9885638, 3.8866415, 3.79134, 3.6935248, 3.5932078, 3.4903867, 3.385059, 3.2775478, 3.1686144, 3.0582895, 2.946573, 2.834149, 2.7226534, 2.612163, 2.502683, 2.3950555, 2.291324, 2.1915886, 2.0958576, 2.004818, 1.9201629, 1.8419797, 1.770277, 1.705355, 1.6479607, 1.5981369, 1.5558903, 1.5210611, 1.4932287, 1.4723767, 1.4585102, 1.451095, 1.448724, 1.4513264, 1.4589053, 1.4707768, 1.4851093, 1.5018047, 1.5208641, 1.541707, 1.5627527, 1.5839117, 1.605183, 1.6262696, 1.6463488, 1.665371, 1.6833333, 1.7002599, 1.7162231, 1.7312256, 1.7452652, 1.7586117, 1.7720442, 1.778811, 1.7924465, 1.8062416, 1.8209932, 1.8370926, 1.854542, 1.8733549, 1.8939221, 1.9164405, 1.9409127, 1.9673413, 1.9957086, 2.0260067, 2.0582385, 2.092402, 2.1283305, 2.1659374, 2.2052233, 2.2461905, 2.2889295, 2.3334875, 2.3798652, 2.4280744, 2.4786181, 2.531767, 2.5875213, 2.645897, 2.707622, 2.773097, 2.8423264, 2.9153225, 2.9924912, 3.0740628, 3.160045, 3.2504346, 3.3446867, 3.4424958, 3.543871, 3.6487937, 3.7554889, 3.8629332, 3.9711378, 4.0800705, 4.187059, 4.290527, 4.3904767, 4.4868703, 4.5770483, 4.659403, 4.733919, 4.806746, 4.8628893, 4.908598, 4.9438477, 4.9686127, 4.982856, 4.9865465, 4.979658, 4.9622254, 4.935879, 4.9013467, 4.8586097, 4.807745, 4.7514243, 4.6908674, 4.6260715, 4.557123, 4.486863, 4.4166255, 4.346408, 4.27628, 4.208481, 4.144081, 4.0830865, 4.0255365, 3.9725912, 3.9248204, 3.8822355, 3.844846, 3.8126547, 3.7856686, 3.763899, 3.7473316, 3.735053, 3.7266092, 3.72201, 3.7212284, 3.722849, 3.7261472, 3.7311277, 3.73776, 3.7446437, 3.751045, 3.7569613, 3.7623744, 3.7662344, 3.7679863, 3.7676265, 3.7651367, 3.7599, 3.7515764, 3.7401586, 3.7256465, 3.7078328, 3.6866047, 3.6619537, 3.6338794, 3.60278, 3.56888, 3.5321944, 3.492728, 3.4515762, 3.4093683, 3.3661058, 3.3218172, 3.2780974, 3.2358787, 3.1951637, 3.15598, 3.1199567, 3.0880666, 3.0603154, 3.0367243, 3.018344, 3.0058138, 2.9991412, 2.9983351, 3.0034857, 3.014652, 3.03184, 3.0550437, 3.0834744, 3.116634, 3.1545281, 3.1971433, 3.2431538, 3.2917078, 3.3428094, 3.3964467, 3.4511683, 3.5060232, 3.561012, 3.616124, 3.6701543, 3.7222977, 3.7725518, 3.8209078, 3.8666832, 3.9094107, 3.9490857, 3.9857018, 4.0191236, 4.0520883, 4.0785975, 4.101815, 4.121998, 4.1392684, 4.153621, 4.1650667, 4.174136, 4.1811075, 4.185973, 4.1887445, 4.190079, 4.1903176, 4.1894593, 4.1875167, 4.185024, 4.1822624, 4.1792336, 4.1759467, 4.172778, 4.169933, 4.1674128, 4.165226, 4.163671, 4.162913, 4.162957, 4.163812, 4.16569, 4.1687055, 4.1728754, 4.1782055, 4.1846786, 4.1923013, 4.201079, 4.211013, 4.221807, 4.233292, 4.245472, 4.2583413, 4.2713923, 4.284323, 4.2907434, 4.303493, 4.3159556, 4.327539, 4.3381863, 4.347891, 4.3565435, 4.363752, 4.369474, 4.3736987, 4.3763857, 4.3774004, 4.3767204, 4.374335, 4.3702946, 4.3648124, 4.357899, 4.34955, 4.3398724, 4.32933, 4.317963, 4.305763, 4.2928696, 4.2798653, 4.2668095, 4.2537017, 4.2406764, 4.228275, 4.2165604, 4.2055383, 4.1952877, 4.186112, 4.1780477, 4.1711035, 4.1652803, 4.1605616, 4.1569514, 4.1544566, 4.1530123, 4.1523294, 4.152378, 4.1531672, 4.154616, 4.156345, 4.158314, 4.160527, 4.1629596, 4.1654906, 4.1681046, 4.1708026, 4.1736646, 4.1770597, 4.1810317, 4.185579, 4.190867, 4.1976657, 4.2060723, 4.2160873, 4.227886, 4.242302, 4.2594433, 4.2793136, 4.3020263, 4.3281083, 4.357637, 4.390617, 4.42704, 4.466849, 4.51004, 4.556618, 4.6064553, 4.6588874, 4.7194595, 4.777163, 4.8370886, 4.89819, 4.9603786, 5.0236573, 5.087708, 5.1513624, 5.214514, 5.2771606, 5.339024, 5.3990736, 5.4572115, 5.513435, 5.5675097, 5.618557, 5.6664906, 5.7113066, 5.7527866, 5.7900996, 5.823157, 5.838087, 5.86474, 5.8865876, 5.903276, 5.914791, 5.92112, 5.9222226, 5.9180665, 5.908636, 5.8939195, 5.8743978, 5.850395, 5.8219013, 5.788913, 5.752312, 5.712712, 5.670105, 5.6244936, 5.5769057, 5.5280685, 5.4779825, 5.426652, 5.3749266, 5.3234234, 5.2721467, 5.221103, 5.1707067, 5.1212645, 5.072781, 5.0252614, 4.97874, 4.933242, 4.8887677, 4.845318, 4.8029017, 4.7615266, 4.721192, 4.6819, 4.643915, 4.6074457, 4.572493, 4.5390606, 4.507611, 4.478514, 4.4517756, 4.4273987, 4.4057064, 4.3869615, 4.3711724, 4.358348, 4.3483987, 4.341247, 4.3368993, 4.335361, 4.3362417, 4.339209, 4.3442674, 4.351419, 4.360289, 4.37055, 4.382203, 4.395248, 4.409571, 4.425072, 4.441751, 4.459607, 4.478773, 4.4993715, 4.5214067, 4.544883, 4.5698833, 4.596487, 4.6247, 4.6545296, 4.685706, 4.717975, 4.7513404, 4.785806, 4.820686, 4.8553185, 4.8897023, 4.923835, 4.943831, 4.9753733, 5.004678, 5.031738, 5.056276, 5.077176, 5.094307, 5.1076574, 5.1171207, 5.1222873, 5.1231017, 5.119552, 5.1117196, 5.099989, 5.0843954, 5.064933, 5.041821, 5.0160384, 4.987697, 4.9567957, 4.923613, 4.8893924, 4.854284, 4.818289, 4.7816577, 4.7455254, 4.7100325, 4.675183, 4.6411314, 4.608588, 4.5776463, 4.5483093, 4.5206146, 4.4947224, 4.4706583, 4.4484262, 4.4279613, 4.4089355, 4.391307, 4.375078, 4.3601427, 4.345964, 4.332469, 4.3196573, 4.3074617, 4.2955446, 4.283859, 4.272403, 4.2611837, 4.250239, 4.239572, 4.229182, 4.219103, 4.2095227, 4.200469, 4.191943, 4.183943, 4.176453, 4.169469, 4.162987, 4.1569595, 4.151133, 4.1454678, 4.139962, 4.1345696, 4.1290326, 4.123313, 4.1174126, 4.111338, 4.1051226, 4.0987706, 4.0922832, 4.085743, 4.079626, 4.074012, 4.0689034, 4.064429, 4.061341, 4.0597677, 4.0597153, 4.0613136, 4.065331, 4.0682974, 4.0761504, 4.0865707, 4.09982, 4.116167, 4.1356163, 4.1581736, 4.1837544, 4.212267, 4.243714, 4.2816954, 4.318839, 4.3581085, 4.3995047, 4.443024, 4.4878354, 4.5333133, 4.579459, 4.626268, 4.67269, 4.7179217, 4.7619596, 4.804797, 4.8454223, 4.883043, 4.917653, 4.9492445, 4.9771194, 5.000721, 5.020041, 5.0350704, 5.045649, 5.0516415, 5.053036, 5.049822, 5.042522, 5.031566, 5.0169425, 4.9986405, 4.9777565, 4.9552226, 4.9310346, 4.9051905, 4.8789496, 4.8534045, 4.828561, 4.8044243, 4.7820587, 4.7623997, 4.745463, 4.7312627, 4.7204776, 4.713719, 4.711001, 4.7123384, 4.71798, 4.728155, 4.742876, 4.7621574, 4.785776, 4.8135214, 4.828944, 4.862896, 4.900842, 4.9419003, 4.9859324, 5.0329432, 5.0827627, 5.1343656, 5.1875825, 5.2424107, 5.2987175, 5.355718, 5.4132843, 5.471416, 5.5300446, 5.5887356, 5.6474195, 5.7061005, 5.7647314, 5.82299, 5.8808265, 5.9382477, 5.995184, 6.05115, 6.1060624, 6.159926, 6.212634, 6.263465, 6.312279, 6.3590665, 6.4037123, 6.4455066, 6.4843035, 6.5200844, 6.552775, 6.581979, 6.607604, 6.6296296, 6.6480494, 6.6629415, 6.6743064, 6.682124, 6.6846967, 6.6875486, 6.687667, 6.685041, 6.6796627, 6.672073, 6.6629333, 6.652245, 6.6400075, 6.6268263, 6.6121016, 6.5985146, 6.5847387, 6.571462, 6.559274, 6.5481796, 6.5381823, 6.529776, 6.5233927, 6.519039, 6.5167203, 6.5165615, 6.518675, 6.5230694, 6.5297537, 6.538412, 6.548754, 6.560787, 6.574515, 6.589325, 6.604644, 6.620474, 6.6368165, 6.6530085, 6.6684203, 6.6830482, 6.69689, 6.7094297, 6.7201695, 6.729106, 6.7362366, 6.741295, 6.744018, 6.7444, 6.7424364, 6.7381454, 6.7315483, 6.722643, 6.7114277, 6.6981707, 6.6831512, 6.66637, 6.647826, 6.627937, 6.607142, 6.585442, 6.562838, 6.539721, 6.516513, 6.493212, 6.469818, 6.4465485, 6.423642, 6.401098, 6.378913, 6.357054, 6.3354855, 6.3142047, 6.2932105, 6.2722325, 6.25096, 6.229389, 6.207519, 6.1849527, 6.1612263, 6.136336, 6.110278, 6.082654, 6.052986, 6.021269, 5.9874973, 5.951425, 5.912749, 5.8714595, 5.8275466, 5.7810884, 5.7321877, 5.680842, 5.627047, 5.5711803, 5.5137224, 5.454673, 5.3940306, 5.332333, 5.2702775, 5.2078686, 5.1451073, 5.0825496, 5.0209293, 4.9602537, 4.9005275, 4.8423085, 4.814045, 4.7592173, 4.706658, 4.656456, 4.6093426, 4.5654902, 4.5249057, 4.487635, 4.45404, 4.424209, 4.3957515, 4.3738356, 4.355619, 4.341096, 4.3302746, 4.323061, 4.31886, 4.3175764, 4.319217, 4.32361, 4.329663, 4.337193, 4.3462048, 4.3564806, 4.366631, 4.376415, 4.385832, 4.394679, 4.4016495, 4.4065056, 4.409241, 4.409738, 4.407259, 4.4016633, 4.392943, 4.3810954, 4.36615, 4.348105, 4.3269544, 4.30279, 4.276283, 4.2475543, 4.2166, 4.1835594, 4.149438, 4.1144314, 4.0785418, 4.0419016, 4.005458, 3.9694002, 3.933731, 3.8985577, 3.864653, 3.8321745, 3.8011246, 3.7716014, 3.7443285, 3.719458, 3.6969953, 3.6770413, 3.660349, 3.6470807, 3.6372426, 3.6309443, 3.629007, 3.631614, 3.6387737, 3.650599, 3.667936, 3.690987, 3.7197735, 3.7543917, 3.7954688, 3.8431451, 3.8974235, 3.9583156, 4.025889, 4.100163, 4.181141, 4.2687244, 4.3620343, 4.460876, 4.5123754, 4.6195383, 4.73119, 4.8458242, 4.96344, 5.0840497, 5.206273, 5.3281083, 5.449546, 5.5705914, 5.6896415, 5.8043294, 5.914633, 6.02055, 6.1205144, 6.212172, 6.295483, 6.370431, 6.435797, 6.4897213, 6.5321493, 6.5630465, 6.5819244, 6.5880375, 6.581335, 6.561773, 6.5298886, 6.48656, 6.4317527, 6.3654222, 6.289121, 6.205403, 6.1142836, 6.0157456, 5.9118505, 5.806024, 5.698327, 5.5887694, 5.4791703, 5.372587, 5.2690864, 5.1588163, 5.0632157, 4.9737616, 4.8904734, 4.8133683, 4.742986, 4.679983, 4.6243773, 4.576183, 4.5352097, 4.5012145, 4.4742103, 4.4542103, 4.440528, 4.432285, 4.429489, 4.43215, 4.43939, 4.450067, 4.464181, 4.481736, 4.5019636, 4.523845, 4.547378, 4.5725646, 4.598885, 4.6256375, 4.652817, 4.6804233, 4.7081757, 4.7356877, 4.7629585, 4.789989, 4.8166647, 4.8428216, 4.8684573, 4.893569, 4.918133, 4.942115, 4.9655156, 4.988336, 5.010538, 5.0320673, 5.0529227, 5.073105, 5.0925393, 5.111116, 5.128831, 5.145683, 5.161638, 5.1766467, 5.190706, 5.203811, 5.216068, 5.227636, 5.2385144, 5.248698, 5.2584662, 5.268261, 5.278087, 5.2879453, 5.2982135, 5.3095016, 5.3218226, 5.3351803, 5.3499627, 5.366804, 5.3857193, 5.406715, 5.4301276, 5.4565167, 5.485898, 5.51828, 5.5538216, 5.5927906, 5.635205, 5.681076, 5.730199, 5.782207, 5.8371086, 5.894917, 5.954995, 6.016201, 6.0785165, 6.1419454, 6.205553, 6.267651, 6.328198, 6.3871846, 6.4436073, 6.49563, 6.5431924, 6.5862746, 6.62403, 6.654895, 6.678802, 6.6957192, 6.705094, 6.705909, 6.69811, 6.681669, 6.656349, 6.617748, 6.5728507, 6.518595, 6.455051, 6.3823256, 6.300405, 6.2092743, 6.1093974, 6.001436, 5.885384, 5.761232, 5.629924, 5.4928308, 5.3499594, 5.2013063, 5.0483117, 4.893098, 4.7356887, 4.576088, 4.4160523, 4.258219, 4.1026244, 3.9492807, 3.7999177, 3.6571767, 3.5211, 3.3917012, 3.2702744, 3.1588311, 3.0574102, 2.966027, 2.885167, 2.8155942, 2.7573352, 2.7104056, 2.6743274, 2.648317, 2.6323764, 2.6265178, 2.629549, 2.639492, 2.6563237, 2.6800504, 2.7093008, 2.7417634, 2.7774048, 2.8162282, 2.8571155, 2.8981464, 2.9392881, 2.98054, 3.021239, 3.0602272, 3.0974815, 3.1329992, 3.1666145, 3.198034, 3.2272491, 3.2542574, 3.2792811, 3.3027265, 3.3246002, 3.3449004, 3.364006, 3.38262, 3.4007583, 3.4184206, 3.4359002, 3.4537475, 3.4719758, 3.490586, 3.5096185, 3.5291514, 3.5391064, 3.5593944, 3.5801504, 3.600855, 3.6213367, 3.6415935, 3.6615462, 3.680054, 3.696737, 3.7115948, 3.7183387, 3.729539, 3.7361357, 3.7380736, 3.735351, 3.726988, 3.7109609, 3.687198, 3.6556888, 3.6157277, 3.560301, 3.499418, 3.4285183, 3.3476813, 3.2570376, 3.156571, 3.0462654, 2.927355, 2.8017566, 2.669488, 2.5305462, 2.3869426, 2.2418478, 2.0953078, 1.9473306, 1.7999429, 1.6563914, 1.5167315, 1.3809743, 1.250666, 1.1884949, 1.0701605, 0.9598435, 0.85765153, 0.7647098, 0.68133503, 0.607532, 0.5432506, 0.4878702, 0.4412166, 0.4032923, 0.38760424, 0.36182395, 0.34217533, 0.32863003, 0.32118833, 0.31889033, 0.32004485, 0.32461995, 0.3326153, 0.34334567, 0.3555816, 0.36225498, 0.37671247, 0.39262944, 0.40972668, 0.42791897, 0.44720665, 0.46765366, 0.4901042, 0.5148219, 0.54180783, 0.57114565, 0.6039605, 0.6406116, 0.681102, 0.72546566, 0.77413297, 0.8272496, 0.8848257, 0.94681215, 1.012328, 1.0810856, 1.1530901, 1.2282138, 1.3044683, 1.381183, 1.4583535, 1.535823, 1.6112534, 1.6838405, 1.753577, 1.8203405, 1.8822882, 1.9387727, 1.9897854, 2.0352683, 2.0743845, 2.1068337, 2.132611, 2.1517282, 2.164471, 2.1709397, 2.17113, 2.1688693, 2.160196, 2.147034, 2.1294267, 2.1073744, 2.081483, 2.0531094, 2.0223053, 1.9890704, 1.9539429, 1.936124, 1.900025, 1.8633127, 1.8260207, 1.7887846, 1.7518517, 1.7152218, 1.678906, 1.64313, 1.6079832, 1.5734657, 1.5564429, 1.5229789, 1.4905189, 1.4590743, 1.4286444, 1.3994389, 1.3719722, 1.3462687, 1.3223284, 1.3110602, 1.2907823, 1.2801197, 1.2648563, 1.2527298, 1.2440555, 1.2394041, 1.2387905, 1.2422173, 1.2495604, 1.2605873, 1.2752961, 1.2936893, 1.3151118, 1.3383293, 1.3633155, 1.3900728, 1.4176328, 1.4441358, 1.4695354, 1.4938306, 1.5161314, 1.5347011, 1.5494925, 1.5605035, 1.5672373, 1.5687071, 1.564881, 1.5557538, 1.5414311, 1.5221307, 1.4978538, 1.4685947, 1.4521976, 1.4172777, 1.3796433, 1.3392924, 1.296324, 1.2523803, 1.2080401, 1.1633054, 1.1182243, 1.0735844, 1.0296688, 0.98647827, 0.944004, 0.9020746, 0.8606265, 0.81965894, 0.7791546, 0.73881257, 0.69852006, 0.6582763, 0.61809605, 0.57826316, 0.5388865, 0.49996784, 0.4615162, 0.42366955, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 2.1568418, 2.2172499, 2.2774363, 2.3370702, 2.3961425, 2.4546473, 2.5126858, 2.570308, 2.6275215, 2.6843686, 2.7416425, 2.7996821, 2.8584971, 2.918117, 2.979055, 3.0415356, 3.1055682, 3.171152, 3.238049, 3.3061566, 3.3754807, 3.4459922, 3.5167553, 3.5873528, 3.657786, 3.7280118, 3.796777, 3.8635092, 3.9282055, 3.9908245, 4.0502343, 4.1059036, 4.1578217, 4.205954, 4.2496095, 4.288456, 4.3224835, 4.3516755, 4.3758087, 4.3947697, 4.4085455, 4.417133, 4.4195714, 4.4208827, 4.41743, 4.409205, 4.3964376, 4.379833, 4.359436, 4.3352427, 4.3075337, 4.2771697, 4.244208, 4.208647, 4.170759, 4.1313896, 4.0905957, 4.048378, 4.0049973, 3.9612799, 3.9172845, 3.873008, 3.8287282, 3.8069155, 3.764015, 3.7220843, 3.6811366, 3.641603, 3.6037235, 3.5675063, 3.532957, 3.5000167, 3.4686506, 3.438861, 3.4106445, 3.383723, 3.3579383, 3.3332906, 3.3097749, 3.287111, 3.2651358, 3.2438476, 3.2232409, 3.2030778, 3.1832192, 3.1636665, 3.1444168, 3.1252384, 3.1059914, 3.086676, 3.0672896, 3.047695, 3.0278063, 3.0055883, 2.9850817, 2.964333, 2.9433641, 2.9221733, 2.9007664, 2.879332, 2.8579562, 2.8366387, 2.8153856, 2.7943685, 2.773668, 2.7532861, 2.73323, 2.7136724, 2.6946929, 2.6762912, 2.6584806, 2.6416645, 2.6260355, 2.6115937, 2.5983636, 2.5924602, 2.5824745, 2.5749192, 2.5697975, 2.5673993, 2.5685763, 2.573388, 2.581838, 2.5941093, 2.6107473, 2.6317935, 2.6572533, 2.6871207, 2.721366, 2.7599921, 2.8030055, 2.8501778, 2.900785, 2.9547803, 3.0121698, 3.0725236, 3.1344593, 3.1978793, 3.2627888, 3.3286464, 3.3936837, 3.4577663, 3.520896, 3.5825744, 3.6411512, 3.6964939, 3.7485998, 3.7734175, 3.8195755, 3.8608294, 3.8971696, 3.9285831, 3.954938, 3.9761517, 3.9922116, 4.0031195, 4.006904, 4.011645, 4.012603, 4.0097666, 4.0036087, 3.9958467, 3.9866283, 3.9759498, 3.964402, 3.9541392, 3.9453607, 3.9415286, 3.9350042, 3.931659, 3.932529, 3.9376233, 3.9469588, 3.9612265, 3.9808693, 4.0059013, 4.0363345, 4.0718827, 4.0915074, 4.1344676, 4.18239, 4.2349687, 4.2909565, 4.350244, 4.4128513, 4.4783697, 4.545104, 4.619722, 4.6886663, 4.758084, 4.8262644, 4.893078, 4.958499, 5.022072, 5.082519, 5.1397424, 5.193725, 5.2443104, 5.291067, 5.312996, 5.3539476, 5.3910227, 5.4245477, 5.4546866, 5.4814353, 5.504806, 5.5254774, 5.5438027, 5.5597825, 5.573435, 5.579604, 5.5909967, 5.6011243, 5.609984, 5.6177406, 5.6249347, 5.6316047, 5.637749, 5.6435266, 5.649457, 5.655583, 5.658719, 5.665153, 5.6724286, 5.680893, 5.690543, 5.701387, 5.7141447, 5.72923, 5.746648, 5.7664084, 5.777273, 5.8011756, 5.827985, 5.8577113, 5.89012, 5.924355, 5.9603534, 5.998129, 6.0371194, 6.075265, 6.1123867, 6.1484914, 6.1829076, 6.21316, 6.2390285, 6.260523, 6.2771406, 6.2869716, 6.289813, 6.28564, 6.2743025, 6.2657638, 6.2428675, 6.212167, 6.173621, 6.1282034, 6.0765476, 6.018629, 5.954444, 5.88584, 5.814045, 5.739055, 5.6608853, 5.581327, 5.5015945, 5.421699, 5.341659, 5.262599, 5.1852913, 5.1097445, 5.0359697, 4.964353, 4.895167, 4.828416, 4.7641034, 4.7020955, 4.642296, 4.5847063, 4.529328, 4.4756813, 4.4234195, 4.372544, 4.347626, 4.298615, 4.2498, 4.20107, 4.1524262, 4.103682, 4.0539756, 4.003202, 3.951363, 3.898378, 3.8713179, 3.8160138, 3.7591288, 3.7006624, 3.6410837, 3.580763, 3.5197005, 3.4578993, 3.3964658, 3.3362913, 3.2715588, 3.2140684, 3.159314, 3.1081274, 3.0605178, 3.016511, 2.9771433, 2.943023, 2.9141583, 2.890562, 2.8724942, 2.8655925, 2.8560586, 2.8522246, 2.853956, 2.86074, 2.8725357, 2.8893497, 2.91098, 2.936656, 2.9663064, 2.9999328, 3.0182316, 3.0573723, 3.0997717, 3.145436, 3.1943686, 3.24629, 3.3010247, 3.3585825, 3.4189672, 3.481624, 3.5461907, 3.5791926, 3.646638, 3.7157476, 3.7854736, 3.855707, 3.9264479, 3.9974241, 4.067526, 4.1366286, 4.204726, 4.271506, 4.3039403, 4.3667526, 4.426817, 4.484118, 4.5378385, 4.587399, 4.632791, 4.674002, 4.710429, 4.741635, 4.767609, 4.7786317, 4.796647, 4.8089013, 4.81533, 4.8159184, 4.810737, 4.8001623, 4.784226, 4.762911, 4.7364845, 4.706231, 4.6723013, 4.634687, 4.5937896, 4.551523, 4.508133, 4.4636207, 4.4183717, 4.374216, 4.3314037, 4.289944, 4.2500534, 4.212736, 4.1781387, 4.1462746, 4.1171575, 4.090802, 4.0672183, 4.0464153, 4.028265, 4.01208, 4.004689, 3.9913127, 3.97981, 3.9695904, 3.9601386, 3.95145, 3.9435194, 3.935925, 3.928295, 3.9198546, 3.9121296, 3.9040196, 3.895315, 3.8860128, 3.8761067, 3.8653502, 3.8535872, 3.8408167, 3.827037, 3.8121707, 3.80431, 3.7877324, 3.770009, 3.7512116, 3.7316353, 3.711309, 3.6902313, 3.66855, 3.6468642, 3.6252382, 3.6036737, 3.5823407, 3.5619345, 3.5425289, 3.5241227, 3.5068676, 3.4914036, 3.477807, 3.4660833, 3.4562864, 3.4486308, 3.4456167, 3.441219, 3.4389987, 3.4386272, 3.439867, 3.4427242, 3.4472003, 3.4525187, 3.4581015, 3.4639494, 3.4669733, 3.472944, 3.4776459, 3.480923, 3.482773, 3.483042, 3.481021, 3.4766161, 3.4698215, 3.460674, 3.4493663, 3.4359162, 3.4283853, 3.4117086, 3.3936987, 3.3750167, 3.355662, 3.3356366, 3.3158972, 3.297231, 3.2796395, 3.2631264, 3.2485592, 3.2366652, 3.2274475, 3.2209103, 3.217631, 3.218107, 3.222346, 3.2303557, 3.2422326, 3.2580605, 3.267458, 3.2892253, 3.3148484, 3.3437297, 3.375786, 3.4110227, 3.4492216, 3.4891713, 3.5306914, 3.573786, 3.6181228, 3.661832, 3.683343, 3.725677, 3.767094, 3.8064585, 3.84269, 3.8757792, 3.9057178, 3.9320033, 3.9541492, 3.972148, 3.9859908, 3.995708, 4.001327, 4.0028386, 4.000232, 3.9939144, 3.9842992, 3.9713826, 3.9551609, 3.9362295, 3.923866, 3.9015856, 3.8772109, 3.850959, 3.823768, 3.7957406, 3.7668715, 3.737414, 3.7085018, 3.6802683, 3.666406, 3.6391933, 3.613491, 3.589924, 3.5684984, 3.54922, 3.5323575, 3.5181172, 3.5065048, 3.4975257, 3.490913, 3.48646, 3.4841716, 3.4840508, 3.4854023, 3.4876738, 3.490869, 3.4949899, 3.4991956, 3.5028002, 3.5058033, 3.5070791, 3.5090044, 3.5092866, 3.507806, 3.5045598, 3.499542, 3.492732, 3.4841223, 3.473708, 3.461599, 3.4483893, 3.4341667, 3.4189348, 3.402814, 3.3864272, 3.369874, 3.3531635, 3.3363683, 3.3198547, 3.3035967, 3.2876546, 3.2720518, 3.25708, 3.2427776, 3.2291365, 3.2162216, 3.204436, 3.1938438, 3.1844451, 3.1762908, 3.169672, 3.1646395, 3.1611977, 3.1600747, 3.1586237, 3.1579742, 3.1581292, 3.159092}
range =
  {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
qp =
  {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
qt =
  {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
qrh =
  {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
qu =
  {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
qv =
  {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
qwind =
  {-999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0}
mr =
  {12.97112, -999.0, -999.0, -999.0, -999.0, -999.0, 12.458791, 12.41971, 12.380868, 12.342213, 12.30434, 12.267463, 12.230986, 12.195017, 12.159777, 12.125516, 12.092484, 12.060945, 12.031214, 12.003624, 11.978735, 11.957224, 11.938713, 11.923472, 11.911771, 11.903867, 11.89997, 11.900279, 11.904986, 11.914232, 11.927921, 11.945893, 11.967984, 11.993983, 12.0234785, 12.056004, 12.091094, 12.128933, 12.168465, 12.208801, 12.249271, 12.289201, 12.327876, 12.364579, 12.398602, 12.4293375, 12.456639, 12.480489, 12.500869, 12.517747, 12.531032, 12.54061, 12.546368, 12.548168, 12.545782, 12.538944, -999.0, 12.5109005, 12.489648, 12.463889, 12.430655, 12.39617, 12.357474, 12.314331, 12.266486, 12.214365, 12.15813, 12.096703, 12.029874, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 10.873554, -999.0, -999.0, -999.0, 10.379188, 10.255982, 10.132407, 10.010559, 9.890429, 9.770604, 9.653895, 9.538589, -999.0, -999.0, -999.0, -999.0, -999.0, 8.899104, 8.804152, 8.714868, 8.62838, 8.54453, 8.464577, 8.387739, -999.0, 8.23961, 8.170104, 8.102508, 8.036688, 7.972688, 7.912335, 7.853901, 7.797252, 7.742403, -999.0, -999.0, 7.5937104, 7.548543, 7.505563, 7.4653196, 7.4281573, 7.3932476, 7.3605595, 7.33004, 7.301633, 7.275266, 7.2510676, 7.2291293, 7.2086906, 7.189595, 7.1717515, 7.1550856, 7.1395254, 7.125026, 7.111696, 7.099687, 7.089155, 7.080235, 7.0729675, 7.0673614, 7.0634255, 7.061234, 7.060537, 7.0610785, 7.062656, 7.065051, 7.067968, 7.071085, 7.0740824, 7.0766463, 7.0784945, 7.0793552, 7.078958, 7.0770965, 7.073908, 7.0696473, 7.0645695, 7.0589194, 7.0529046, 7.046096, 7.039939, 7.034013, 7.028511, 7.0236287, 7.01956, 7.0164814, 7.0144997, 7.013702, 7.0141745, 7.015949, 7.0188246, 7.0225396, 7.0268316, 7.031433, 7.0360394, 7.040337, 7.0440154, 7.0467973, 7.0485473, 7.049168, 7.0485644, 7.0466537, 7.043418, 7.038856, 7.0329666, 7.025734, 7.0170765, 7.006895, 6.995088, 6.981621, 6.9667673, 6.9508934, 6.9349647, 6.918767, 6.9026628, 6.887025, 6.872226, 6.858591, 6.846212, 6.835112, 6.825314, 6.8167596, 6.8089886, 6.8014193, 6.7934713, 6.78462, 6.7745967, 6.7634263, 6.750989, 6.736917, 6.7213497, 6.7045126, 6.6866317, 6.6679163, 6.6484976, 6.628483, 6.607979, 6.587081, 6.5658183, 6.544906, 6.523635, 6.502015, 6.4801025, 6.457969, 6.435688, 6.413329, 6.3909583, 6.3686395, 6.3468323, 6.325552, 6.3045216, 6.283818, 6.263519, 6.2436633, 6.2240667, 6.2044625, 6.184582, 6.1641603, 6.1434894, 6.122038, 6.099393, 6.0753865, 6.050182, 6.0240645, 5.9973245, 5.970274, 5.943907, 5.9184537, 5.8940597, 5.8711658, 5.8499947, 5.830687, 5.8133807, 5.798189, 5.785072, 5.773928, 5.7647657, 5.7575464, 5.7520323, 5.7482333, 5.746156, 5.745848, 5.7476006, 5.7523675, 5.7596955, 5.770259, 5.7844734, 5.803066, 5.826032, 5.853655, 5.886024, 5.9231644, 5.96509, 6.012041, 6.0648346, 6.122031, 6.1833506, 6.249188, 6.319797, 6.3933554, 6.4698367, -999.0, -999.0, 6.7160683, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 6.650762, 6.6113124, 6.5738187, 6.5386257, 6.5029597, 6.473687, 6.448166, 6.4257216, 6.406451, 6.3902087, 6.376763, 6.365877, 6.3573065, 6.3507776, 6.346007, 6.342715, -999.0, -999.0, 6.338404, 6.3375072, 6.336237, 6.3343215, -999.0, -999.0, -999.0, -999.0, 6.3082895, 6.2988734, 6.287799, 6.2751617, 6.2611146, 6.245809, 6.229405, 6.212115, 6.1941733, 6.175814, 6.157256, 6.139201, 6.1212783, 6.103464, 6.0858665, 6.068689, 6.0521727, 6.036559, 6.022097, 6.0090785, 5.997812, 5.9886055, 5.981752, 5.9774427, 5.9759526, 5.977227, 5.981393, 5.9885454, 5.998889, 6.012342, 6.028912, 6.04847, 6.0708327, 6.0958138, 6.123204, 6.1526494, 6.183738, 6.2160625, 6.249718, 6.2844477, 6.3195367, 6.3547564, 6.3898773, 6.424646, 6.4588013, 6.49248, 6.5255766, 6.5573177, 6.587522, 6.6160116, 6.6426272, 6.6673417, 6.690183, 6.711177, 6.7303576, 6.7479124, 6.764213, 6.779036, 6.792537, 6.805005, 6.816784, 6.8282127, 6.8395944, 6.8510194, 6.862483, 6.873985, 6.8855286, 6.89715, 6.9089036, 6.92085, -999.0, -999.0, 6.959981, 6.9736304, 6.9879427, 7.0028872, 7.01839, 7.0343795, 7.050744, 7.0671515, 7.083193, 7.0984635, 7.112618, 7.1256237, 7.1375623, 7.1485105, 7.158615, 7.167996, 7.1767693, 7.1851063, 7.193174, 7.201146, 7.209197, 7.2174973, 7.2262, 7.2353544, 7.24497, 7.2550545, 7.2656054, 7.2765493, 7.287787, 7.2992196, 7.310724, 7.3220143, -999.0, -999.0, 7.3511796, 7.3583107, 7.3637543, 7.367298, 7.368759, 7.3681393, 7.365515, 7.3609624, 7.354567, 7.346495, 7.3369474, 7.326553, 7.315195, 7.3030596, 7.290435, 7.277606, 7.2648497, 7.252376, 7.2403655, 7.2289987, 7.2184362, 7.208704, 7.1997695, 7.1915994, 7.1841583, 7.1773944, 7.171247, 7.1659737, 7.161199, 7.156781, 7.1525774, 7.1484485, 7.1442637, 7.139963, 7.1355166, 7.130895, 7.1260767, 7.121086, 7.1159697, 7.110773, 7.105524, 7.1000934, 7.094281, 7.0878906, 7.080715, 7.0724645, 7.0628095, 7.051421, 7.038289, 7.0231752, 7.005527, 6.985075, -999.0, -999.0, 6.905017, 6.871925, -999.0, -999.0, -999.0, -999.0, -999.0, 6.6159143, 6.5648203, -999.0, -999.0, 6.3955007, 6.3358946, 6.2744145, -999.0, -999.0, 6.0874586, -999.0, 5.9665294, 5.9097624, 5.855236, 5.8035197, 5.7522893, 5.7096295, 5.6709347, 5.6364837, 5.606777, 5.582113, 5.561461, 5.544582, 5.5312114, 5.5210023, 5.513565, 5.5085063, -999.0, -999.0, -999.0, 5.5053115, 5.5074124, 5.5101876, 5.513431, 5.51694, 5.5205274, 5.5240993, 5.527602, 5.530986, 5.5342307, 5.5375404, 5.5412173, 5.54556, 5.5508647, 5.5574193, 5.565505, 5.5754, 5.5873537, 5.601433, 5.617619, 5.6358933, 5.656199, 5.6782093, 5.701474, 5.7258344, 5.751029, 5.776204, 5.800962, 5.824913, 5.8476934, 5.8691115, -999.0, -999.0, -999.0, 5.9389863, 5.9521165, 5.963566, 5.972998, 5.9806004, 5.986672, 5.99151, 5.9953995, 5.9985533, 6.0011473, 6.0033555, 6.005331, 6.0070505, 6.008402, 6.009272, -999.0, -999.0, 6.0081944, 6.0065107, 6.004141, 6.0011587, 5.997735, 5.9940934, 5.9901876, 5.9860125, 5.981508, 5.9766126, 5.9712586, 5.965302, 5.95856, -999.0, 5.942011, 5.9320774, 5.92119, 5.909491, 5.8971257, 5.8842783, 5.8711543, 5.8579583, 5.8448925, 5.832425, 5.8205934, 5.8093514, 5.797833, 5.7882037, 5.779405, 5.7714643, 5.7643886, 5.758045, 5.7522397, 5.746778, 5.741482, 5.736277, 5.7311373, 5.726036, 5.7209554, 5.7159333, 5.7110343, 5.7063227, 5.7018566, 5.6976466, 5.6936803, 5.6899467, 5.6864815, 5.6833773, 5.6804857, 5.677807, 5.6753454, 5.673161, 5.671339, 5.669966, 5.6691155, 5.6687584, 5.668816, 5.669214, 5.669874, 5.670703, 5.6715965, 5.672453, 5.6731644, 5.6735888, 5.673565, 5.67293, 5.6715336, 5.6693316, 5.6663313, 5.662541, 5.6579633, 5.652564, 5.64629, 5.639087, 5.6309223, 5.621926, 5.6123176, 5.6023164, 5.592135, 5.5819244, 5.572188, 5.5627003, 5.5535226, 5.544701, 5.5362487, 5.5281787, 5.520517, 5.5134053, 5.5070477, 5.501648, 5.497412, 5.4945645, 5.493339, 5.4939694, 5.496663, 5.501394, 5.5080013, 5.5163207, 5.5261865, 5.537435, 5.549904, 5.56343, 5.5778513, 5.5930414, 5.608896, 5.6253147, 5.642211, 5.6595984, 5.6775494, 5.69629, 5.7160974, 5.736574, 5.757585, 5.7789936, 5.800645, 5.822165, 5.8430495, 5.8627963, 5.8809314, 5.897246, 5.9116926, 5.9242277, 5.934811, 5.9434624, 5.95024, 5.9552, 5.958401, 5.9599285, 5.9598, 5.9581494, 5.9551563, 5.9510274, 5.9460173, 5.9403806, 5.934369, 5.9282193, 5.92216, 5.91642, 5.911215, 5.9066486, 5.902767, 5.8996167, 5.8972354, 5.895598, 5.894646, 5.8943214, 5.8945613, 5.8952756, 5.8963594, 5.897708, 5.899217, 5.900792, 5.9023423, 5.9037766, 5.9050026, 5.9058967, 5.906319, 5.90613, 5.9051957, 5.903443, 5.9008303, 5.8973165, 5.8928666, 5.8875237, 5.8813705, 5.8744917, 5.86697, 5.8588758, 5.850274, 5.8412285, 5.831807, 5.8220954, 5.8124976, 5.8028607, 5.79323, 5.78371, 5.7744083, 5.7654343, 5.7568917, 5.748827, 5.744978, 5.7376523, 5.7308326, 5.7245107, 5.7186327, 5.71314, 5.7079725, 5.703066, 5.698346, 5.693738, 5.6891656, 5.684594, 5.6800804, 5.675695, 5.671509, 5.6675906, 5.6640034, 5.6608105, 5.658074, 5.6558127, 5.653941, 5.652358, 5.650982, 5.6497917, 5.64868, 5.6476274, 5.6466146, 5.64561, 5.6445546, 5.643384, 5.642036, 5.6404324, 5.6384616, 5.636006, -999.0, -999.0, 5.6248083, 5.61977, 5.614127, 5.607935, 5.601318, 5.5944104, 5.587347, 5.5802693, 5.5733376, 5.566714, 5.5605617, 5.555013, 5.550118, 5.545913, 5.542128, 5.539458, 5.537456, 5.5360494, 5.5351663, 5.534707, 5.5345197, 5.534555, 5.534556, 5.534369, 5.5338683, 5.5329313, 5.531435, 5.5292897, -999.0, -999.0, 5.5188165, 5.5139484, 5.508386, 5.5021296, 5.4951797, 5.487485, 5.478879, 5.469179, 5.4582024, 5.4457865, 5.4318137, 5.416171, 5.398746, 5.380097, 5.3596144, 5.3371973, 5.3127894, 5.28633, 5.2577577, 5.2270055, 5.194793, 5.160712, 5.1243815, 5.085785, 5.0449004, 5.0029073, 4.9590573, -999.0, 4.8651285, 4.816725, 4.766894, 4.7156844, -999.0, -999.0, 4.560895, 4.5090756, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 4.1800966, 4.1409674, 4.104192, 4.070048, 4.039059, 4.0115504, 3.9868991, 3.9651334, 3.946127, 3.9297218, 3.9157543, 3.9041843, 3.8948374, 3.8871658, 3.880914, 3.8758118, 3.8715546, 3.867832, 3.8643332, 3.8607664, 3.8568876, 3.8524609, -999.0, -999.0, -999.0, 3.825635, 3.8163285, 3.8059664, 3.7946663, 3.782656, 3.7703776, 3.7576, 3.7444894, 3.7312162, 3.7179532, 3.7048779, 3.6921828, 3.6800632, 3.6687155, 3.658322, 3.6493883, 3.6416583, 3.635247, 3.6302812, 3.6266382, 3.6251125, 3.6254115, 3.6275883, 3.6315517, 3.6371896, -999.0, 3.652984, 3.6627061, 3.6732712, 3.6843994, 3.6960704, -999.0, -999.0, 3.7307317, 3.7413294, 3.7512138, 3.7603016, 3.7685113, 3.7757332, 3.78179, 3.7864964, 3.7896695, 3.7911656, 3.790933, 3.7889318, 3.7851222, 3.7794805, -999.0, -999.0, 3.7518249, 3.739143, 3.725042, 3.7099373, 3.6935666, 3.6760612, 3.6575649, 3.6382248, 3.6181874, 3.5977108, 3.5776396, 3.5675776, 3.547557, 3.5278785, 3.508671, -999.0, -999.0, -999.0, 3.4388795, 3.4232366, 3.4081614, 3.3936386, 3.3796751, 3.3662958, 3.3535833, -999.0, -999.0, 3.3205514, 3.310827, 3.301762, 3.2933834, 3.285729, 3.2788377, 3.2727454, 3.2674541, 3.2629378, 3.259167, 3.2561057, 3.2536597, 3.2516913, 3.2501736, 3.2488425, -999.0, 3.2461255, 3.2444193, 3.2422698, 3.2395217, 3.2360246, 3.2316287, -999.0, 3.2196805, 3.212154, 3.2036698, 3.1942887, 3.184113, 3.1732793, 3.1619246, 3.150345, 3.138749, 3.1268299, 3.1145818, 3.1019974, 3.0890515, 3.075706, 3.061921, 3.0476553, 3.0333345, 3.0185547, 3.0031674, 2.9871233, 2.970401, 2.953004, 2.934986, 2.9169621, -999.0, -999.0, -999.0, 2.839887, 2.8202698, 2.8011181, 2.7822373, 2.7638419, 2.7461276, 2.727641, 2.7124932, 2.6985917, 2.6859915, 2.6747606, 2.664963, 2.6566556, 2.6498325, 2.6444414, 2.6404266, 2.637727, 2.636253, 2.635947, 2.6365807, 2.6380355, 2.6401975, 2.642955, 2.6461985, 2.6498275, 2.653813, 2.6580257, 2.6601946, 2.664613, 2.66909, 2.6735973, 2.6781127, 2.682614, 2.6870792, 2.691483, 2.6958013, 2.7000096, 2.7040768, 2.70795, 2.7115734, 2.7148917, 2.7178578, 2.7204475, 2.7226408, 2.7244182, 2.7257671, 2.726695, 2.7272136, 2.7273335, 2.7270696, 2.726446, 2.7254891, 2.7242248, 2.722688, 2.720944, 2.7190633, 2.7171156, 2.7151783, 2.7133722, 2.7118773, 2.710689, 2.7099097, 2.7096498, 2.7100217, 2.7111363, 2.7130785, 2.7158515, 2.7194421, 2.7238362, 2.7289977, 2.7348561, 2.7413826, 2.748333, -999.0, -999.0, -999.0, 2.7793322, 2.7879028, 2.7968428, 2.8061867, 2.8159685, 2.826202, 2.8368335, 2.8477962, 2.859024, 2.870448, 2.882343, 2.8942597, 2.9061089, 2.9178076, 2.9292924, 2.9405053, 2.9513893, 2.9619205, 2.9721928, 2.9823248, 2.9924335, 3.0026278, 3.013066, 3.0240028, 3.035276, 3.0469313, 3.0588894, 3.0710433, 3.083287, 3.0954988, 3.1074924, 3.119068, 3.1300275, 3.1362314, 3.1458905, 3.1546507, 3.1625242, 3.1694984, 3.1754727, 3.1805563, 3.184858, 3.1884885, 3.1915846, 3.1943052, 3.1968083, 3.199246, -999.0, -999.0, -999.0, 3.2096152, 3.2125375, 3.2156348, 3.218921, 3.2224107, 3.226113, 3.2300334, 3.2341778, 3.2385523, 3.243162, 3.2480109, 3.2531033, 3.2584398, 3.2639666, 3.2695854, 3.2751975, 3.2807047, 3.2860045, 3.2909887, 3.2955508, 3.2995872, 3.3030438, 3.305909, 3.3081713, 3.309821, 3.3108835, 3.3114152, 3.311473, 3.3111134, 3.3104033, 3.3094187, 3.3082347, 3.306926, 3.3055477, 3.304137, 3.3027303, 3.301363, 3.3000395, 3.2987382, 3.2974348, 3.2961059, 3.2947142, 3.2932122, 3.2915509, 3.2896833, 3.28759, 3.2852786, 3.2827568, 3.2800345, 3.2772224, 3.274424, 3.2716167, 3.2688737, 3.2662926, 3.2639935, 3.2620976, 3.2607229, 3.2599354, 3.2597501, 3.26018, 3.261236, 3.262896, 3.2651067, 3.2678125, 3.2709596, 3.2744944, 3.2763903, 3.2804067, 3.284679, 3.2891526, 3.2937653, 3.2984514, 3.303146, 3.3077846, 3.312303, 3.316637, 3.3211143, 3.324855, 3.3282313, 3.3311975, 3.3337228, 3.3357396, 3.3372235, 3.338193, 3.3386276, 3.3385127, 3.3378475, 3.3366323, 3.334868, 3.3325496, 3.3296556, 3.3261614, 3.322042, 3.317264, 3.311767, 3.3054838, 3.298348, 3.290286, 3.2812026, 3.2709973, 3.2595692, 3.2468169, 3.233166, 3.2180986, 3.2014642, 3.1831717, 3.163161, 3.1413765, 3.1182437, 3.093744, 3.0675662, 3.0398483, -999.0, 2.9816658, 2.9515553, 2.9208465, 2.8902717, 2.8604686, 2.8309634, 2.802029, 2.774593, 2.7486422, 2.7239847, 2.7008302, 2.679647, 2.6608653, 2.6439643, 2.6362267, 2.6221912, 2.6100903, 2.5998707, 2.5914083, 2.5847828, 2.5797017, 2.575945, 2.5733984, 2.5719469, 2.5714765, 2.5719135, 2.573225, 2.5753794, 2.5783455, 2.5821085, 2.586671, 2.5920362, 2.5982072, 2.6051917, 2.6130018, 2.6216958, 2.6314738, 2.6421115, 2.6535547, 2.6657472, 2.678632, 2.69209, 2.705936, 2.7199833, 2.7340481, 2.7479506, 2.7617471, 2.775198, 2.7879374, 2.79982, 2.8107347, 2.8205729, 2.8292255, 2.8366168, 2.842707, 2.8474572, 2.8493176, 2.851997, 2.8533266, 2.8533607, 2.8521528, 2.8497624, 2.8462787, 2.8417995, 2.8364232, 2.8302464, 2.8226383, 2.815081, 2.8070474, 2.7989364, 2.790459, 2.7816584, 2.7725787, 2.7632582, 2.7537146, 2.7439609, 2.7340097, 2.7238705, 2.7136905, 2.7036152, 2.6933322, 2.682831, 2.6720982, 2.6611202, 2.6498833, 2.6383767, 2.6266053, 2.6150582, 2.603308, 2.591325, 2.5791175, 2.566694, 2.5540626, 2.5412335, 2.52853, 2.5159192, 2.5031705, 2.4903004, 2.4773207, 2.4642408, 2.451071, 2.4382112, 2.425469, 2.4126813, 2.3998644, 2.387043, 2.3742807, 2.361651, 2.349723, 2.3380997, 2.3268027, 2.3158884, 2.3054137, 2.2954278, 2.2859435, 2.2770486, 2.2689643, 2.2613654, 2.25421, 2.2474456, 2.2410197, 2.2348778, 2.228955, 2.2231834, 2.217495, 2.211827, 2.206141, 2.200651, 2.1951168, 2.189478, 2.1837332, 2.1778889, 2.17195, 2.1659229, 2.1598105, 2.1536155, 2.147341, 2.1409912, 2.1345773, 2.1284094, 2.122211, 2.1159885, 2.1097567, 2.1035314, 2.097328, 2.0911605, 2.085036, 2.0789597, 2.0729363, 2.0669708, 2.0611804, 2.0556185, 2.0501263, 2.0447092, 2.039375, 2.034132, 2.028989, 2.023953, 2.021474, 2.0165904, 2.0118005, 2.0070975, 2.0024712, 1.9979064, 1.993447, 1.9891726, 1.9849175, 1.980678, 1.9760289, 1.9718121, 1.9675997, 1.9633857, 1.9591638, 1.9549279, 1.9506732, 1.9463964, 1.9420941, 1.9377632, 1.9334047, 1.9290239, 1.9247835, 1.9205813, 1.9163629, 1.912113, 1.907816, 1.9034566, 1.8990221, 1.8945034, 1.8898909, 1.8851757, 1.8803527, 1.8754209, 1.8703793, 1.8652272, 1.8600746, 1.8549402, 1.84969, 1.8443202, 1.838828, 1.833211, 1.8274667, 1.8215932, 1.8155886, 1.8094524, 1.8031842, 1.796783, 1.790477, 1.7841134, 1.777636, 1.7710514, 1.7643727, 1.7576214, 1.7508192, 1.743988, 1.7371472, 1.7303134, 1.7236942, 1.7172146, 1.7107909, 1.7044427, 1.6981897, 1.6920518, 1.6860517, 1.6802162, 1.674572, 1.6691471, 1.6640031, 1.6594094, 1.6553341, 1.6518277, 1.6489049, 1.6464785, 1.6444551, 1.6427407, 1.6412423, 1.6398679, 1.6385252, 1.6371226, 1.6355932, 1.6339006, 1.6329827, 1.6309819, 1.628735, 1.6262211, 1.6234235, 1.620325, 1.6169118, 1.6131862, 1.6092281, 1.6051164, 1.6007298, 1.5960815, 1.5911866, 1.58606, 1.5807166, 1.575172, 1.5694418, 1.5635419, 1.5574886, 1.5514668, 1.5454636, 1.5393709, 1.5332079, 1.5269916, 1.5207376, 1.5144621, 1.5081804, 1.5019014, 1.4958318, 1.4898782, 1.4839475, 1.4780542, 1.4722152, 1.4664472, 1.4607668, 1.4551864, 1.4497168, 1.4444414, 1.4394705, 1.4346232, 1.4298942, 1.4248223, 1.420324, 1.4159287, 1.411633, 1.4074332, 1.4033254, 1.3993051, 1.3953671, 1.3916023, 1.3879958, 1.3844504, 1.3809578, 1.3775095, 1.3740966, 1.3707095, 1.3673376, 1.3639702, 1.3605977, 1.3572134, 1.3538119, 1.3503873, 1.3469352, 1.3434781, 1.3401396, 1.3367741, 1.3333818, 1.3299648, 1.326525, 1.3230649, 1.319587, 1.3160958, 1.3125962, 1.3090931, 1.3055906, 1.302087, 1.2985786, 1.2951217, 1.2917686, 1.2883918, 1.2849783, 1.2815142, 1.2779869, 1.274387, 1.2707068, 1.2669381, 1.2630737, 1.2591109, 1.2550484, 1.2508851, 1.2467674, 1.2426134, 1.2383671, 1.2340316, 1.2296101, 1.2251074, 1.2205285, 1.2158788, 1.2111628, 1.2063808, 1.2016059, 1.1969208, 1.1921703, 1.1873581, 1.1824894, 1.1775688, 1.1726013, 1.1675922, 1.1625457, 1.157467, 1.1525944, 1.1477212, 1.1428548, 1.1380129, 1.1332154, 1.128496, 1.123894, 1.1194487, 1.1151998, 1.1112863, 1.1077349, 1.1044881, 1.1015816, 1.09903, 1.09684, 1.0950179, 1.0935645, 1.0924462, 1.091615, 1.091023, 1.090621, 1.0903547, 1.0901673, 1.0900023, 1.0898033, 1.0895157, 1.0890856, 1.088459, 1.0875851, 1.0864315, 1.0849742, 1.0832312, 1.0812259, 1.0786322, 1.0759302, 1.0729083, 1.0695765, 1.0659575, 1.0620779, 1.0579644, 1.0536449, 1.0491513, 1.0445585, 1.0400447, 1.0354601, 1.0308379, 1.0262108, 1.021612, 1.0170735, 1.0126209, 1.0082777, 1.0040953, 1.0002337, 0.99653, 0.9929922, 0.9896281, 0.9864429, 0.9834284, 0.9805717, 0.97785956, 0.9752774, 0.972802, 0.9704069, 0.9680655, 0.9657519, 0.9635184, 0.9613016, 0.95904756, 0.9567354, 0.95434433, 0.9518536, 0.9492423, 0.94649154, 0.94359505, 0.94055116, 0.93735826, 0.93401647, 0.93053734, 0.926937, 0.9233326, 0.91971236, 0.91601676, 0.9122545, 0.9084344, 0.9045663, 0.90066665, 0.89675456, 0.8928492, 0.8889698, 0.8852112, 0.88161635, 0.87810415, 0.8746925, 0.87138915, 0.8681976, 0.8651216, 0.86216307, 0.85931313, 0.8565586, 0.8538862, 0.8512822, 0.8488126, 0.8464179, 0.84403914, 0.8416597, 0.83926463, 0.83805674, 0.8356114, 0.8331148, 0.8305596, 0.82794994, 0.82529074, 0.8225872, 0.81984496, 0.81707054, 0.8143646, 0.81302536, 0.8103361, 0.8076342, 0.80492055, 0.80219615, 0.79946244, 0.79672444, 0.793989, 0.7912629, 0.7885537, 0.7856073, 0.7829827, 0.7805332, 0.7781531, 0.7758591, 0.7736687, 0.7715995, 0.7696681, 0.76788443, 0.7662562, 0.76479113, 0.7634944, 0.76235735, 0.7613662, 0.76050717, 0.7597647, 0.7591129, 0.7585223, 0.75796324, 0.7574061, 0.7571192, 0.7565108, 0.7558323, 0.7550548, 0.7541503, 0.7530922, 0.751854, 0.7504674, 0.748868, 0.7470396, 0.744972, 0.7438452, 0.7414025, 0.73872095, 0.735821, 0.7327234, 0.72945064, 0.72603416, 0.7225092, 0.71891105, 0.71534204, 0.71186584, 0.7101397, 0.7067345, 0.703423, 0.70023763, 0.6972035, 0.6943451, 0.6916866, 0.68924606, 0.6870321, 0.6850523, 0.68332547, 0.6819, 0.6807119, 0.6797619, 0.6790509, 0.67859095, 0.67841154, 0.67854387, 0.67901856, 0.67982894, 0.6809078, 0.68218213, 0.68357897, 0.68504965, 0.6865238, 0.6878872, 0.6890599, 0.6899906, 0.69067526, 0.6911148, 0.6913103, 0.69127214, 0.69102675, 0.6906019, 0.6900256, 0.6893273, 0.6885393, 0.68769413, 0.68684137, 0.68602246, 0.68523127, 0.6844905, 0.6841461, 0.6835225, 0.6829951, 0.68257236, 0.6822631, 0.68207526, 0.68201256, 0.6820766, 0.68226886, 0.68259096, 0.6828008, 0.68331796, 0.68396485, 0.68474126, 0.6856434, 0.6866611, 0.68778354, 0.68899995, -999.0, -999.0, -999.0, -999.0, 0.69561076, 0.6972906, 0.69902194, 0.7007956, 0.70260274, 0.7044394, 0.70630413, 0.7081953, 0.7091504, 0.71107894, 0.7122479, 0.71421576, 0.7162081, 0.7182237, 0.72025377, 0.72228646, 0.7243099, 0.7263116, 0.7282758, 0.7302636, 0.73217756, 0.7339991, 0.7357241, 0.7373537, 0.7388891, 0.7403318, 0.7416873, 0.7429624, 0.74416393, 0.7452986, 0.7463721, 0.7473894, 0.74835557, 0.74927664, 0.75016373, 0.7510305, 0.75189054, 0.7527578, 0.7536491, 0.7545824, 0.75557566, 0.7561003, 0.75721276, 0.75841385, 0.7597091, 0.76110387, 0.76259875, 0.7641858, 0.7658563, 0.7676016, 0.7694194, 0.7713416, 0.773279, 0.7752068, 0.7770983, 0.778924, 0.78065383, 0.7822579, 0.7837117, 0.7850002, 0.78610975, 0.7870265, 0.7877471, 0.788287, 0.7886637, 0.78889483, 0.7890069, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 0.8829371, 0.8830745, 0.8828777, 0.88230354, 0.8813113, 0.8798602, 0.87794894, 0.87565297, 0.87305695, 0.8702456, 0.86728954, 0.86423117, 0.86110955, 0.85796374, 0.85482526, 0.8517503, 0.8488173, 0.8459339, 0.8431088, 0.84034, 0.83762443, 0.83495885, 0.83233964, 0.8297621, 0.82722133, 0.82471246, 0.82222986, 0.8197666, 0.81734157, 0.8150166, 0.8126896, 0.8103527, 0.80799806, 0.8056179, 0.80320436, 0.8007492, 0.7982441, 0.7956809, 0.793052, 0.79035145, 0.7875732, 0.78475654, 0.7833663, 0.7805276, 0.7776175, 0.77464384, 0.77161425, 0.7685373, 0.7654219, 0.76227707, 0.7591115, 0.7559315, 0.75278056, 0.7497418, 0.7467023, 0.74366707, 0.7406415, 0.737631, 0.7346408, 0.73167086, 0.72871864, 0.72578126, 0.72285634, 0.72143775, 0.71867734, 0.7159386, 0.7132268, 0.7105476, 0.7079084, 0.7053165, 0.70277935, 0.70030296, 0.69789, 0.6955424, 0.69326234, 0.69109565, 0.6890564, 0.6870775, 0.6851565, 0.6832896, 0.6814709, 0.67969376, 0.6779518, 0.6762396, 0.6745539, 0.6728918, 0.67125064, 0.669629, 0.668029, 0.6664536, 0.66490555, 0.6634094, 0.6620011, 0.6604892, 0.6591506, 0.65784603, 0.6565716, 0.65532297, 0.65409565, 0.6528854, 0.6516884, 0.65050083, 0.64931893, 0.64814013, 0.6469643, 0.6457919, 0.64462304, 0.6434582, 0.64229757, 0.6411416, 0.6399905, 0.6388452, 0.6377077, 0.6366305, 0.6355742, 0.63505095, 0.6340134, 0.6329864, 0.6319683, 0.63095737, 0.6299513, 0.6289477, 0.6279439, 0.62693715, 0.6259221, 0.6248916, 0.62383854, 0.622756, 0.62163824, 0.62048054, 0.619278, 0.6180261, 0.6167238, 0.61537224, 0.61397254, 0.6125259, 0.61108303, 0.60962546, 0.60812795, -999.0, -999.0, 0.6034354, 0.6018314, 0.60022205, 0.5986134, 0.59700954, 0.5954147, 0.59462196, 0.5930471, 0.5914855, -999.0, -999.0, -999.0, -999.0, -999.0, 0.5825429, 0.58181053, 0.58032966, 0.5788186, 0.5772673, 0.5756657, 0.5740087, 0.5722944, 0.5705212, 0.5686873, 0.56679326, 0.56484085, 0.56384337, 0.5618886, 0.5599044, 0.5578647, 0.55576634, 0.5536056, 0.55138224, 0.5491042, 0.546781, 0.54442203, 0.542039, 0.5408438, 0.5384906, 0.5362431, 0.53403425, 0.53188777, 0.52983093, 0.5278914, 0.52609575, 0.5244567, -999.0, 0.52153254, 0.52038705, 0.5193645, 0.51840895, 0.51746416, 0.5165219, 0.51552767, 0.51445395, 0.513289, 0.51202184, 0.5106501, 0.50992584, 0.5084023, 0.506781, 0.5050675, 0.5032739, 0.50141317, 0.4994983, 0.49754015, 0.49561766, 0.49369493, 0.491745, 0.49076086, 0.48877373, 0.48675984, 0.48471728, 0.48264417, 0.48053938, 0.4784023, 0.47623223, 0.47414696, 0.47202918, 0.4698765, 0.46878657, 0.46657854, 0.4643318, 0.4620455, 0.45971885, 0.45735115, 0.45499256, 0.45266265, 0.45028502, 0.447856, 0.4466212, 0.44410998, 0.44154224, 0.43891674, 0.4362324, 0.4336212, 0.43097234, 0.4282776, 0.42554134, 0.4227717, 0.41997948, 0.41717562, 0.41448852, 0.41185063, 0.40926442, 0.40675962, 0.4043649, 0.40209332, 0.39994672, 0.397955, 0.39616743, 0.39531547, 0.39368024, 0.39211634, 0.39059937, 0.38911036, 0.38764575, 0.38620475, 0.38478658, 0.3833905, 0.38201633, 0.3807385, 0.37947965, 0.37823987, 0.37702087, 0.3758247, 0.3746535, 0.37350872, 0.37239042, 0.37129834, 0.3702322, 0.36919087, 0.368171, 0.3671687, 0.36619085, 0.3652702, 0.36435395, 0.36343727, 0.36251542, 0.3615831, 0.36063355, 0.3596596, 0.3591613, 0.3581376, 0.35707477, 0.35597068, 0.35482332, 0.3536309, 0.35239476, 0.35111892, 0.34986705, 0.3485946, 0.34794882, 0.34664246, 0.34532225, 0.34399527, 0.3426685, 0.3413487, 0.34004265, 0.33875707, 0.33749807, 0.33626965, 0.33497015, 0.33387956, 0.3328277, 0.33181587, 0.33084524, 0.32991692, 0.32903162, 0.3281889, 0.3273882, 0.32662883, 0.3259095, 0.32556373, 0.32489762, 0.3242622, 0.32365355, 0.32306826, 0.32250315, 0.32195503, 0.32142088, 0.32089964, 0.3203993, 0.3199345, 0.31970716, 0.31926295, 0.31883344, 0.3184194, 0.31802166, 0.31764132, 0.31728023, 0.31694028, 0.31662348, 0.31633142, 0.31606454, 0.31594062, 0.31571212, 0.31550932, 0.3153289, 0.31516504, 0.3150118, 0.31486306, 0.3147108, 0.31454536, 0.31435713, 0.3141366, 0.31401196, 0.31373128, 0.31340492, 0.31302842, 0.31259876, 0.31211713, 0.31158543, 0.31100568, 0.3103796, 0.30970812, 0.3090211, 0.30866995, 0.30793676, 0.30716234, 0.3063462, 0.30548787, 0.3045868, 0.30364242, 0.30265403, 0.3016209, 0.30054238, 0.299419, 0.29825208, 0.29704309, 0.29581955, 0.29460412, 0.29335812, 0.29208636, 0.29079387, 0.28948635, 0.28817022, 0.2868519, 0.28553793, 0.28423518, 0.2829511, 0.28174472, 0.28058583, 0.2794652, 0.2783888, 0.27736256, 0.27639225, 0.27548015, 0.27504563, 0.27421907, 0.27344823, 0.27273113, 0.27206233, 0.27143565, 0.27084485, 0.27028376, 0.26976946, 0.26923507, 0.26876116, 0.26829308, 0.26782596, 0.26735497, 0.2668753, 0.26638308, 0.26587713, 0.2653566, 0.2648208, 0.2642696, 0.26398867, 0.26341742, 0.26283517, 0.26224384, 0.26164448, 0.26103762, 0.26042372, 0.2598032, 0.2591755, 0.2585605, 0.25795257, 0.2573337, 0.25670266, 0.2560584, 0.25539973, 0.25472566, 0.2540367, 0.25333446, 0.25262067, 0.25189704, 0.25116578, 0.25079814, 0.25006038, 0.2493216, 0.248584, 0.24784851, 0.24712546, 0.24643703, 0.24575303, 0.24507648, 0.2444107, 0.24408288, 0.24343944, 0.24281332, 0.24220486, 0.24161428, 0.24104181, 0.24048644, 0.2399462, 0.23941907, 0.23890305, 0.23839577, 0.23789461, 0.23764549, -999.0, 0.23665133, 0.23616803, 0.23569441, 0.23521586, 0.23473123, 0.23424053, 0.23374408, 0.23324214, 0.232735, 0.23222281, 0.2317058, 0.23118412, 0.23065785, 0.23012646, 0.22958937, 0.229046, 0.22849591, 0.22793947, 0.22765903, 0.22709402, 0.22652392, 0.22594902, 0.22540182, 0.224853, 0.22429991, 0.22374249, 0.22318052, 0.22261375, -999.0, 0.22146593, 0.22117665, 0.22059646, 0.22001524, 0.21943389, 0.2188516, 0.21826714, 0.2176793, 0.21708721, 0.21649101, 0.21589121, 0.21532184, 0.21475297, 0.21418194, -999.0, -999.0, -999.0, -999.0, 0.21130067, 0.21071571, 0.2101257, 0.20976895, 0.2091694, 0.20856307, 0.2079493, 0.20732671, 0.20669338, 0.20605507, 0.2054319, 0.20479275, 0.20413554, 0.20379949, 0.20311114, 0.2024, 0.20166637, 0.20091096, 0.20013446, 0.19933783, 0.1985228, 0.19769135, 0.19684535, 0.19600745, 0.19518535, 0.1943519, 0.19350739, 0.19265246, -999.0, -999.0, -999.0, -999.0, -999.0, 0.1873907, 0.18694866, 0.18610273, 0.18527262, -999.0, -999.0, -999.0, 0.1820744, 0.18132481, -999.0, -999.0, 0.17925704, 0.178638, 0.17805767, 0.17752801, 0.17706363, 0.17664793, 0.17628685, 0.17598593, -999.0, 0.17554778, 0.1753907, 0.17526163, 0.17515223, 0.1750558, 0.17496571, 0.17487542, 0.17478134, 0.17468256, 0.17457837, 0.17446806, 0.17435202, 0.17423163, 0.17410839, 0.17404613, 0.17392105, 0.1737954, 0.1736693, 0.17354287}
vt =
  {303.75998, -999.0, -999.0, -999.0, -999.0, -999.0, 303.7783, 303.74042, 303.7015, 303.6614, 303.62003, 303.57727, 303.53302, 303.48727, 303.44003, 303.39142, 303.34152, 303.2905, 303.2386, 303.1862, 303.13358, 303.08115, 303.0291, 302.97778, 302.92746, 302.87836, 302.83066, 302.7846, 302.74033, 302.698, 302.65753, 302.61884, 302.58185, 302.54642, 302.51242, 302.4797, 302.4481, 302.41748, 302.38776, 302.35876, 302.33047, 302.30276, 302.2755, 302.24863, 302.22202, 302.1956, 302.1694, 302.14352, 302.118, 302.09296, 302.06842, 302.0446, 302.02148, 301.9993, 301.97815, 301.95828, -999.0, 301.9231, 301.90833, 301.89587, 301.88525, 301.87878, 301.8756, 301.87598, 301.8801, 301.88824, 301.90045, 301.91672, 301.9371, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 302.37283, -999.0, -999.0, -999.0, 302.50925, 302.54025, 302.56934, 302.5957, 302.61844, 302.63684, 302.6507, 302.6598, -999.0, -999.0, -999.0, -999.0, -999.0, 302.6186, 302.5988, 302.5759, 302.55, 302.5212, 302.48972, 302.45578, -999.0, 302.38132, 302.34116, 302.29913, 302.2553, 302.2098, 302.16263, 302.11374, 302.0632, 302.011, -999.0, -999.0, 301.8463, 301.78937, 301.7317, 301.67334, 301.61444, 301.55518, 301.4957, 301.43634, 301.37738, 301.3191, 301.26175, 301.2057, 301.1512, 301.0986, 301.04803, 300.99966, 300.95367, 300.91016, 300.8691, 300.83057, 300.7944, 300.76062, 300.729, 300.6993, 300.6713, 300.64468, 300.6193, 300.5948, 300.57095, 300.5475, 300.52423, 300.50092, 300.47733, 300.4533, 300.42877, 300.4036, 300.37778, 300.35126, 300.32404, 300.29608, 300.26743, 300.23813, 300.2082, 300.1746, 300.14355, 300.11212, 300.08035, 300.04846, 300.0165, 299.98465, 299.95294, 299.9215, 299.89035, 299.85956, 299.82904, 299.79874, 299.76855, 299.73837, 299.70813, 299.67773, 299.64713, 299.6162, 299.58493, 299.5532, 299.521, 299.48822, 299.45477, 299.42047, 299.3852, 299.3488, 299.31113, 299.27203, 299.23132, 299.18893, 299.1448, 299.099, 299.05154, 299.00253, 298.95215, 298.90063, 298.84827, 298.79526, 298.74207, 298.68912, 298.63687, 298.5858, 298.53598, 298.48758, 298.44073, 298.3955, 298.35208, 298.31058, 298.27112, 298.2338, 298.1986, 298.16537, 298.134, 298.10434, 298.07617, 298.04926, 298.0234, 297.99832, 297.9739, 297.95, 297.92657, 297.90347, 297.8808, 297.8586, 297.83704, 297.81616, 297.796, 297.77658, 297.75784, 297.7398, 297.72232, 297.7052, 297.6883, 297.6714, 297.65436, 297.637, 297.6192, 297.60083, 297.58173, 297.5619, 297.5412, 297.51965, 297.49728, 297.47418, 297.45044, 297.4262, 297.4015, 297.3764, 297.351, 297.32535, 297.2995, 297.27353, 297.24747, 297.22147, 297.1955, 297.16968, 297.14404, 297.11868, 297.09363, 297.0689, 297.04462, 297.02072, 296.99738, 296.97238, 296.95047, 296.92938, 296.9092, 296.89005, 296.87198, 296.85507, 296.83932, 296.82477, 296.8113, 296.799, 296.78775, 296.7775, 296.76813, 296.75964, 296.75195, 296.74512, 296.7391, -999.0, -999.0, 296.72617, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 296.31583, 296.27856, 296.23944, 296.1982, 296.1502, 296.10394, 296.0551, 296.00354, 295.94916, 295.8922, 295.83292, 295.7716, 295.70856, 295.64404, 295.57843, 295.512, -999.0, -999.0, 295.3101, 295.24237, 295.17465, 295.1072, -999.0, -999.0, -999.0, -999.0, 294.78473, 294.7242, 294.6651, 294.60718, 294.55026, 294.4941, 294.4385, 294.3832, 294.32803, 294.27277, 294.21725, 294.1614, 294.10526, 294.0488, 293.99207, 293.9353, 293.8789, 293.82315, 293.76843, 293.71518, 293.66388, 293.615, 293.569, 293.52603, 293.48624, 293.44968, 293.4164, 293.38644, 293.35965, 293.336, 293.3153, 293.29733, 293.28156, 293.2676, 293.25504, 293.24335, 293.23212, 293.2208, 293.20895, 293.1963, 293.1826, 293.16766, 293.15128, 293.13324, 293.11337, 293.09146, 293.06732, 293.04074, 293.01157, 292.97958, 292.9446, 292.9065, 292.86508, 292.82022, 292.7718, 292.7197, 292.66388, 292.60434, 292.54095, 292.4739, 292.40326, 292.32913, 292.2517, 292.17123, 292.088, 292.00235, 291.91455, 291.8252, 291.73502, 291.64465, -999.0, -999.0, 291.37, 291.2848, 291.20197, 291.12155, 291.0435, 290.96768, 290.89407, 290.82248, 290.75262, 290.68433, 290.61737, 290.55164, 290.487, 290.42343, 290.3608, 290.2991, 290.2382, 290.17804, 290.11856, 290.05972, 290.00146, 289.94373, 289.88647, 289.82962, 289.773, 289.7166, 289.66028, 289.60394, 289.54752, 289.49097, 289.43414, 289.37704, -999.0, -999.0, 289.20325, 289.14426, 289.08463, 289.02423, 288.96307, 288.90103, 288.83817, 288.7744, 288.70978, 288.64432, 288.57803, 288.511, 288.44327, 288.37488, 288.306, 288.23666, 288.16702, 288.09717, 288.0272, 287.9572, 287.8874, 287.81772, 287.74826, 287.67902, 287.61005, 287.54132, 287.47278, 287.40442, 287.33618, 287.26804, 287.20004, 287.13214, 287.06436, 286.99673, 286.92926, 286.862, 286.79498, 286.72827, 286.66193, 286.59604, 286.53064, 286.4659, 286.40207, 286.33926, 286.27774, 286.21774, 286.1596, 286.10364, 286.05017, 285.99942, 285.95166, 285.90707, -999.0, -999.0, 285.79437, 285.76416, -999.0, -999.0, -999.0, -999.0, -999.0, 285.65833, 285.65082, -999.0, -999.0, 285.6341, 285.62836, 285.62152, -999.0, -999.0, 285.58932, -999.0, 285.55524, 285.5339, 285.50986, 285.48325, 285.45114, 285.41968, 285.3864, 285.35162, 285.31564, 285.27866, 285.2408, 285.20224, 285.16302, 285.12317, 285.08255, 285.0411, -999.0, -999.0, -999.0, 284.86575, 284.81958, 284.77258, 284.7249, 284.6767, 284.62808, 284.57925, 284.53033, 284.4815, 284.43295, 284.3849, 284.3376, 284.29123, 284.24606, 284.20227, 284.16, 284.1194, 284.08054, 284.04352, 284.00836, 283.975, 283.94354, 283.9138, 283.88565, 283.85892, 283.83347, 283.80914, 283.7857, 283.76297, 283.74072, 283.71884, -999.0, -999.0, -999.0, 283.632, 283.60974, 283.58707, 283.56378, 283.53986, 283.51526, 283.48996, 283.4639, 283.4371, 283.40952, 283.3812, 283.35208, 283.32217, 283.29138, 283.2597, -999.0, -999.0, 283.1586, 283.12268, 283.0855, 283.04712, 283.00748, 282.96658, 282.92447, 282.88116, 282.8367, 282.7911, 282.74448, 282.6968, 282.6482, -999.0, 282.54837, 282.49734, 282.44565, 282.39346, 282.34088, 282.28802, 282.23502, 282.18207, 282.12927, 282.07675, 282.0245, 281.9726, 281.91592, 281.86484, 281.81424, 281.7642, 281.71472, 281.66577, 281.61734, 281.56937, 281.52176, 281.47452, 281.4276, 281.381, 281.33475, 281.2888, 281.24313, 281.19778, 281.1527, 281.10785, 281.06296, 281.01797, 280.97263, 280.92676, 280.88013, 280.83252, 280.7837, 280.73383, 280.68323, 280.6322, 280.58105, 280.53006, 280.47943, 280.42947, 280.3804, 280.33224, 280.28488, 280.23828, 280.19232, 280.1467, 280.10104, 280.05493, 280.008, 279.96002, 279.91083, 279.8603, 279.8082, 279.75452, 279.6991, 279.64188, 279.5828, 279.52213, 279.4602, 279.3975, 279.33432, 279.27112, 279.20828, 279.1462, 279.0853, 279.02582, 278.968, 278.91202, 278.85815, 278.80655, 278.75745, 278.711, 278.66736, 278.62668, 278.58893, 278.55423, 278.5225, 278.49332, 278.46594, 278.43967, 278.41376, 278.38776, 278.36127, 278.33395, 278.30548, 278.276, 278.24585, 278.21545, 278.18518, 278.15546, 278.12668, 278.09924, 278.07358, 278.0497, 278.02753, 278.0069, 277.9877, 277.96957, 277.95215, 277.93497, 277.9176, 277.89993, 277.88193, 277.86362, 277.84497, 277.82605, 277.8069, 277.78757, 277.76807, 277.74857, 277.72714, 277.7079, 277.6889, 277.67026, 277.65195, 277.63403, 277.6165, 277.5994, 277.58276, 277.5667, 277.55124, 277.53638, 277.5222, 277.5087, 277.49588, 277.48373, 277.47217, 277.46112, 277.45047, 277.44022, 277.4303, 277.42065, 277.41125, 277.4021, 277.39322, 277.3846, 277.3763, 277.36832, 277.3606, 277.3532, 277.34607, 277.33923, 277.33264, 277.32635, 277.32028, 277.31448, 277.30887, 277.30347, 277.29825, 277.29312, 277.28806, 277.28302, 277.27792, 277.2727, 277.26733, 277.26172, 277.2558, 277.24948, 277.24274, 277.23547, 277.22763, 277.2192, 277.2148, 277.20563, 277.19595, 277.18588, 277.1754, 277.1646, 277.1535, 277.14215, 277.13055, 277.11868, 277.10657, 277.09418, 277.08154, 277.0686, 277.0554, 277.04187, 277.02795, 277.01364, 276.99884, 276.9835, 276.96753, 276.95087, 276.93344, 276.9152, 276.89603, 276.87595, 276.8549, 276.8328, 276.80975, 276.7858, 276.761, 276.73538, 276.70895, 276.68173, -999.0, -999.0, 276.59534, 276.56506, 276.53415, 276.5026, 276.4705, 276.43796, 276.40506, 276.37186, 276.3385, 276.30502, 276.27158, 276.23822, 276.20508, 276.1722, 276.13654, 276.10464, 276.0734, 276.04288, 276.01324, 275.9846, 275.95706, 275.93076, 275.90582, 275.8824, 275.86053, 275.84045, 275.82224, 275.80594, -999.0, -999.0, 275.76776, 275.75818, 275.74966, 275.74176, 275.73413, 275.72626, 275.7178, 275.70834, 275.6974, 275.68466, 275.66998, 275.65314, 275.634, 275.61252, 275.58875, 275.5628, 275.53485, 275.50507, 275.47357, 275.44064, 275.4065, 275.3713, 275.33536, 275.29892, 275.2622, 275.22552, 275.18893, -999.0, 275.11667, 275.08118, 275.04623, 275.01178, -999.0, -999.0, 274.91144, 274.87833, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 274.62897, 274.58984, 274.55023, 274.5103, 274.47037, 274.4306, 274.39133, 274.35275, 274.31494, 274.27798, 274.24203, 274.2071, 274.17316, 274.14017, 274.1081, 274.07687, 274.04633, 274.0163, 273.98663, 273.95715, 273.92767, 273.89813, -999.0, -999.0, -999.0, 273.7765, 273.74493, 273.71283, 273.68018, 273.647, 273.61328, 273.57907, 273.54434, 273.50903, 273.47318, 273.43677, 273.39984, 273.36252, 273.32486, 273.28696, 273.2489, 273.21085, 273.17285, 273.13504, 273.09357, 273.05594, 273.01834, 272.98065, 272.94287, 272.9049, -999.0, 272.82837, 272.7897, 272.7508, 272.7116, 272.67215, -999.0, -999.0, 272.55112, 272.50964, 272.46765, 272.42508, 272.38205, 272.33862, 272.29492, 272.2511, 272.20734, 272.16382, 272.12082, 272.07867, 272.0377, 271.99814, -999.0, -999.0, 271.89014, 271.85837, 271.82898, 271.8021, 271.77786, 271.75635, 271.73767, 271.72192, 271.70917, 271.6995, 271.69296, 271.6909, 271.68912, 271.6906, 271.69522, -999.0, -999.0, -999.0, 271.7403, 271.7569, 271.77505, 271.79446, 271.81476, 271.83563, 271.8568, -999.0, -999.0, 271.9183, 271.93658, 271.95297, 271.96698, 271.97824, 271.98633, 271.99088, 271.9917, 271.98877, 271.9821, 271.97165, 271.95755, 271.94, 271.91922, 271.89532, -999.0, 271.8393, 271.80762, 271.77386, 271.73828, 271.70108, 271.66254, -999.0, 271.58234, 271.5413, 271.50003, 271.45886, 271.41806, 271.37796, 271.33878, 271.3008, 271.26425, 271.22922, 271.19583, 271.1642, 271.13437, 271.10626, 271.07983, 271.05505, 271.03177, 271.00983, 270.98898, 270.96912, 270.95004, 270.93158, 270.91367, 270.89612, -999.0, -999.0, -999.0, 270.82596, 270.80737, 270.78796, 270.7674, 270.74548, 270.72205, 270.69446, 270.66757, 270.63898, 270.60864, 270.57663, 270.54294, 270.5077, 270.47092, 270.43274, 270.39328, 270.35263, 270.31094, 270.26828, 270.2248, 270.18057, 270.13574, 270.09033, 270.0444, 269.99802, 269.9512, 269.904, 269.88025, 269.8325, 269.78442, 269.73605, 269.68744, 269.63864, 269.58963, 269.5405, 269.49124, 269.44193, 269.39255, 269.34314, 269.29373, 269.24435, 269.19504, 269.14584, 269.09686, 269.04813, 268.99976, 268.95178, 268.9042, 268.85715, 268.81058, 268.76453, 268.71896, 268.6739, 268.62927, 268.58508, 268.54123, 268.49768, 268.45438, 268.41132, 268.36844, 268.3257, 268.28314, 268.24078, 268.19873, 268.157, 268.11572, 268.0749, 268.0346, 267.9949, 267.95584, 267.91736, 267.8794, 267.8419, -999.0, -999.0, -999.0, 267.6952, 267.65897, 267.62283, 267.58682, 267.5509, 267.5151, 267.47943, 267.4439, 267.40848, 267.37323, 267.33813, 267.30313, 267.26828, 267.23352, 267.1989, 267.16443, 267.1301, 267.09598, 267.0621, 267.02853, 266.99536, 266.96265, 266.93042, 266.89877, 266.86777, 266.83737, 266.80756, 266.77817, 266.74915, 266.7203, 266.6915, 266.66245, 266.63293, 266.6149, 266.58423, 266.55267, 266.52014, 266.48648, 266.45172, 266.4158, 266.37885, 266.3408, 266.30176, 266.26172, 266.2207, 266.1788, -999.0, -999.0, -999.0, 266.00415, 265.95947, 265.9148, 265.87033, 265.8263, 265.7829, 265.74026, 265.69855, 265.65787, 265.61832, 265.5799, 265.54254, 265.50632, 265.4712, 265.43716, 265.40417, 265.37228, 265.3414, 265.31155, 265.2827, 265.25482, 265.22784, 265.2017, 265.17633, 265.1516, 265.1276, 265.10422, 265.0815, 265.0595, 265.03827, 265.01788, 264.99838, 264.97995, 264.96252, 264.9461, 264.93066, 264.9161, 264.90237, 264.88925, 264.87656, 264.86407, 264.85156, 264.8387, 264.82516, 264.8106, 264.79483, 264.77768, 264.759, 264.73868, 264.71674, 264.69336, 264.66864, 264.64282, 264.61603, 264.58847, 264.56036, 264.53186, 264.50314, 264.4744, 264.4457, 264.41724, 264.3892, 264.3617, 264.3349, 264.30905, 264.2842, 264.27225, 264.24918, 264.2274, 264.207, 264.18793, 264.1701, 264.15347, 264.13788, 264.12317, 264.1091, 264.09402, 264.08044, 264.06665, 264.05243, 264.0374, 264.0214, 264.00418, 263.9856, 263.96545, 263.94366, 263.9201, 263.89478, 263.8676, 263.83862, 263.80783, 263.7753, 263.7411, 263.70526, 263.6679, 263.6291, 263.5889, 263.5474, 263.5046, 263.46057, 263.41534, 263.36896, 263.32135, 263.2725, 263.2224, 263.171, 263.1181, 263.06363, 263.00735, 262.9492, 262.88922, 262.8275, -999.0, 262.69952, 262.63376, 262.56735, 262.50076, 262.4344, 262.36865, 262.30396, 262.2407, 262.17926, 262.1199, 262.06284, 262.00836, 261.9566, 261.90756, 261.884, 261.8388, 261.79605, 261.75552, 261.71692, 261.67996, 261.6443, 261.60965, 261.5759, 261.54282, 261.51025, 261.47806, 261.44635, 261.4151, 261.38434, 261.35422, 261.32483, 261.2964, 261.269, 261.2429, 261.21823, 261.19522, 261.17407, 261.15488, 261.13773, 261.12265, 261.10968, 261.09872, 261.08957, 261.08197, 261.07574, 261.0706, 261.06622, 261.06235, 261.05865, 261.05487, 261.0507, 261.0458, 261.03995, 261.03284, 261.02426, 261.014, 261.00818, 260.995, 260.9798, 260.96255, 260.94333, 260.9221, 260.899, 260.8741, 260.84763, 260.8196, 260.78717, 260.75632, 260.72427, 260.69113, 260.6569, 260.62164, 260.58533, 260.54803, 260.5097, 260.47037, 260.42993, 260.38843, 260.34576, 260.30188, 260.25668, 260.2101, 260.16214, 260.1128, 260.06204, 260.0099, 259.95636, 259.9015, 259.8453, 259.78784, 259.72916, 259.66928, 259.60828, 259.5462, 259.48315, 259.4192, 259.35443, 259.28897, 259.2229, 259.1564, 259.0895, 259.02243, 258.95526, 258.8882, 258.82144, 258.75516, 258.6896, 258.62503, 258.56168, 258.49982, 258.43954, 258.38092, 258.3241, 258.26907, 258.21585, 258.1643, 258.1144, 258.06607, 258.01913, 257.97342, 257.9288, 257.88507, 257.84207, 257.79962, 257.75757, 257.71573, 257.674, 257.6324, 257.59082, 257.54926, 257.50763, 257.466, 257.42432, 257.3826, 257.34076, 257.29874, 257.2565, 257.214, 257.17123, 257.12836, 257.08545, 257.04254, 256.99976, 256.9572, 256.915, 256.87326, 256.832, 256.7913, 256.7512, 256.71176, 256.67297, 256.6349, 256.59747, 256.56076, 256.52475, 256.48947, 256.4549, 256.42102, 256.40436, 256.3715, 256.3393, 256.30765, 256.27655, 256.24588, 256.21555, 256.18546, 256.15555, 256.12573, 256.09305, 256.0633, 256.0335, 256.00363, 255.97359, 255.94331, 255.9128, 255.882, 255.85092, 255.81952, 255.78781, 255.7558, 255.72353, 255.69102, 255.65826, 255.62521, 255.59181, 255.558, 255.52379, 255.48921, 255.4543, 255.4191, 255.38362, 255.34792, 255.312, 255.27592, 255.23967, 255.20325, 255.16663, 255.1298, 255.09279, 255.05557, 255.01817, 254.98059, 254.94283, 254.90485, 254.86664, 254.82817, 254.78941, 254.75037, 254.711, 254.6713, 254.63127, 254.59096, 254.5504, 254.50964, 254.46872, 254.42769, 254.38657, 254.34543, 254.3043, 254.26332, 254.22256, 254.18217, 254.14229, 254.10315, 254.06494, 254.02794, 253.99265, 253.95988, 253.93057, 253.90553, 253.8849, 253.86795, 253.85391, 253.84196, 253.83134, 253.82127, 253.81099, 253.79971, 253.78691, 253.77232, 253.7643, 253.74661, 253.72662, 253.7043, 253.67966, 253.65276, 253.62363, 253.59242, 253.55927, 253.5243, 253.48773, 253.44968, 253.41032, 253.36986, 253.32845, 253.28621, 253.24323, 253.19962, 253.15546, 253.11081, 253.06575, 253.02031, 252.97455, 252.92853, 252.8823, 252.83594, 252.78949, 252.74303, 252.6966, 252.65022, 252.60399, 252.55798, 252.51234, 252.46718, 252.4226, 252.37872, 252.33557, 252.29323, 252.25175, 252.2111, 252.17123, 252.1282, 252.0898, 252.05203, 252.0149, 251.9784, 251.94249, 251.90717, 251.87236, 251.83803, 251.80412, 251.77057, 251.73727, 251.70413, 251.67107, 251.63799, 251.60484, 251.57155, 251.53807, 251.50435, 251.47043, 251.4363, 251.40195, 251.36739, 251.33263, 251.29771, 251.2626, 251.22734, 251.19188, 251.15622, 251.12035, 251.0843, 251.04808, 251.01173, 250.97528, 250.93877, 250.90225, 250.86575, 250.82935, 250.793, 250.75671, 250.72047, 250.68427, 250.64809, 250.6119, 250.5757, 250.53949, 250.50323, 250.46692, 250.43051, 250.39401, 250.35738, 250.3206, 250.28365, 250.2465, 250.20918, 250.17168, 250.13402, 250.0962, 250.05823, 250.02008, 249.98175, 249.9432, 249.9045, 249.86562, 249.82663, 249.78755, 249.74847, 249.70952, 249.6708, 249.63243, 249.5945, 249.5571, 249.52032, 249.48428, 249.449, 249.41452, 249.38087, 249.34807, 249.31613, 249.28503, 249.25479, 249.22534, 249.19664, 249.16856, 249.14099, 249.11382, 249.0868, 249.05977, 249.03247, 249.00465, 248.97615, 248.94676, 248.91629, 248.88455, 248.85135, 248.81645, 248.77965, 248.74072, 248.69958, 248.6562, 248.6105, 248.56248, 248.50711, 248.4546, 248.40024, 248.34418, 248.28667, 248.22798, 248.16837, 248.10811, 248.04749, 247.98676, 247.92624, 247.86621, 247.80698, 247.74883, 247.6921, 247.63707, 247.58395, 247.53296, 247.48427, 247.43805, 247.39438, 247.3533, 247.31482, 247.27896, 247.24557, 247.21448, 247.18547, 247.15834, 247.13283, 247.1086, 247.08533, 247.06274, 247.0406, 247.01872, 246.99689, 246.97495, 246.95271, 246.93005, 246.90681, 246.88289, 246.8582, 246.83273, 246.80649, 246.77942, 246.7516, 246.72308, 246.69394, 246.66425, 246.63399, 246.60318, 246.57181, 246.53989, 246.50748, 246.47469, 246.4416, 246.40833, 246.37497, 246.34166, 246.30853, 246.27568, 246.24321, 246.21114, 246.17953, 246.14844, 246.11784, 246.0877, 246.058, 246.02867, 245.99968, 245.97092, 245.9423, 245.91376, 245.88521, 245.8709, 245.84215, 245.81319, 245.78394, 245.75438, 245.72455, 245.69443, 245.664, 245.63322, 245.60208, 245.58636, 245.5546, 245.52245, 245.48996, 245.4572, 245.42424, 245.39117, 245.35808, 245.32506, 245.2922, 245.25645, 245.22443, 245.19301, 245.16234, 245.13261, 245.10402, 245.07675, 245.05098, 245.02689, 245.00461, 244.98431, 244.96614, 244.95016, 244.93645, 244.92502, 244.91594, 244.90909, 244.90433, 244.90152, 244.90048, 244.90056, 244.90169, 244.9039, 244.90686, 244.91026, 244.91371, 244.91681, 244.91917, 244.92038, 244.92, 244.91759, 244.91548, 244.90923, 244.90009, 244.88797, 244.87274, 244.85432, 244.83281, 244.80843, 244.78137, 244.75185, 244.72026, 244.70383, 244.66997, 244.63515, 244.59988, 244.56467, 244.53004, 244.49657, 244.46472, 244.43495, 244.4077, 244.38338, 244.36241, 244.34511, 244.33179, 244.32278, 244.31857, 244.31987, 244.32742, 244.34196, 244.36351, 244.39091, 244.42296, 244.45836, 244.49577, 244.53363, 244.57036, 244.60439, 244.63457, 244.66052, 244.6819, 244.69838, 244.70981, 244.71635, 244.71822, 244.7156, 244.70877, 244.69814, 244.68414, 244.6672, 244.64777, 244.62633, 244.60338, 244.59149, 244.5672, 244.54251, 244.51775, 244.49324, 244.4693, 244.44614, 244.4239, 244.40273, 244.38275, 244.37325, 244.35522, 244.33856, 244.3233, 244.3095, 244.29706, 244.28601, 244.27628, -999.0, -999.0, -999.0, -999.0, 244.24792, 244.24484, 244.24286, 244.24191, 244.24199, 244.24304, 244.24504, 244.24799, 244.24979, 244.25407, 244.25708, 244.26279, 244.26935, 244.27676, 244.28487, 244.2935, 244.30246, 244.31157, 244.32054, 244.32907, 244.33685, 244.34361, 244.34924, 244.35374, 244.35706, 244.35918, 244.3602, 244.3602, 244.35931, 244.35764, 244.35532, 244.3525, 244.34933, 244.34601, 244.34271, 244.3397, 244.33722, 244.3355, 244.33478, 244.33536, 244.33746, 244.33917, 244.344, 244.35074, 244.35947, 244.37022, 244.38298, 244.39757, 244.41382, 244.43152, 244.45045, 244.47028, 244.49062, 244.51115, 244.5315, 244.55124, 244.56995, 244.5872, 244.60268, 244.6162, 244.62758, 244.63667, 244.64346, 244.64813, 244.65096, 244.65216, 244.6521, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 245.70938, 245.70654, 245.69894, 245.68604, 245.66731, 245.64227, 245.61092, 245.57437, 245.53381, 245.4905, 245.4454, 245.39912, 245.35219, 245.30516, 245.25844, 245.21225, 245.1668, 245.12225, 245.07875, 245.03627, 244.99477, 244.95421, 244.91457, 244.87572, 244.83759, 244.80008, 244.76312, 244.72656, 244.69029, 244.65419, 244.61813, 244.58202, 244.54572, 244.50912, 244.47214, 244.43462, 244.39645, 244.35753, 244.31773, 244.27698, 244.2352, 244.19234, 244.17047, 244.12596, 244.0805, 244.03424, 243.98729, 243.93979, 243.8919, 243.84375, 243.7955, 243.74722, 243.699, 243.65092, 243.60303, 243.55539, 243.50806, 243.46104, 243.41443, 243.36823, 243.32243, 243.27707, 243.23215, 243.20987, 243.1657, 243.12207, 243.07907, 243.03673, 242.99512, 242.95428, 242.91426, 242.87514, 242.83698, 242.79984, 242.76382, 242.72897, 242.69527, 242.66267, 242.63115, 242.60066, 242.57112, 242.54239, 242.51439, 242.487, 242.46016, 242.43378, 242.4078, 242.38217, 242.35689, 242.332, 242.3075, 242.28343, 242.25984, 242.2345, 242.21204, 242.19017, 242.16887, 242.14807, 242.12773, 242.10782, 242.08824, 242.0689, 242.04968, 242.03056, 242.01149, 241.99242, 241.97333, 241.95422, 241.93509, 241.91594, 241.89679, 241.87766, 241.8586, 241.83965, 241.82089, 241.81158, 241.79309, 241.77477, 241.75653, 241.73836, 241.7202, 241.70195, 241.68356, 241.66496, 241.64607, 241.6268, 241.60706, 241.58676, 241.56587, 241.54436, 241.5222, 241.49937, 241.47585, 241.45161, 241.42665, 241.40091, 241.3744, 241.34709, 241.31894, -999.0, -999.0, 241.22989, 241.1991, 241.16801, 241.13673, 241.10535, 241.0739, 241.05818, 241.02678, 240.99544, -999.0, -999.0, -999.0, -999.0, -999.0, 240.80826, 240.79253, 240.7608, 240.72864, 240.69583, 240.66225, 240.6278, 240.59245, 240.55617, 240.5189, 240.48068, 240.44153, 240.42162, 240.38113, 240.33978, 240.29749, 240.2541, 240.20955, 240.16376, 240.11688, 240.0691, 240.0206, 239.9716, 239.94702, 239.89793, 239.84924, 239.80133, 239.75467, 239.7098, 239.66727, 239.62761, 239.59108, -999.0, 239.52464, 239.49788, 239.47353, 239.45042, 239.42744, 239.40346, 239.37794, 239.3507, 239.32147, 239.2901, 239.25655, 239.23897, 239.20227, 239.16357, 239.123, 239.08081, 239.0373, 238.9927, 238.9473, 238.90112, 238.85425, 238.80676, 238.7828, 238.73442, 238.6854, 238.63568, 238.5852, 238.53397, 238.48192, 238.42908, 238.37541, 238.3209, 238.26558, 238.23761, 238.18106, 238.12373, 238.06573, 238.00716, 237.94815, 237.88876, 237.82901, 237.7689, 237.7084, 237.67801, 237.61679, 237.55486, 237.49197, 237.42793, 237.3627, 237.2963, 237.22874, 237.1601, 237.09055, 237.02036, 236.94981, 236.87921, 236.80911, 236.74036, 236.67369, 236.60992, 236.54941, 236.49226, 236.43858, 236.38843, 236.3646, 236.31902, 236.27568, 236.23398, 236.19337, 236.1538, 236.11514, 236.07738, 236.04047, 236.00435, 235.96896, 235.93431, 235.90033, 235.86702, 235.83443, 235.80255, 235.7714, 235.74094, 235.71114, 235.68199, 235.65343, 235.62537, 235.59769, 235.57027, 235.54301, 235.5158, 235.4885, 235.46098, 235.43312, 235.40472, 235.3756, 235.3607, 235.33011, 235.2984, 235.26552, 235.23146, 235.19618, 235.15974, 235.12227, 235.0839, 235.04471, 235.02489, 234.9849, 234.94464, 234.90437, 234.86429, 234.82457, 234.78539, 234.74689, 234.70924, 234.67255, 234.63339, 234.59904, 234.56596, 234.53418, 234.50372, 234.47466, 234.44696, 234.42064, 234.39566, 234.37196, 234.34953, 234.33876, 234.31798, 234.29817, 234.27919, 234.26093, 234.24324, 234.22603, 234.20917, 234.19263, 234.17644, 234.16063, 234.15286, 234.13766, 234.12292, 234.10867, 234.09494, 234.08179, 234.06926, 234.0574, 234.04628, 234.03592, 234.02632, 234.02179, 234.01329, 234.0055, 233.99828, 233.99146, 233.98483, 233.97823, 233.97136, 233.96393, 233.95561, 233.9461, 233.94083, 233.92915, 233.91588, 233.90086, 233.88403, 233.8654, 233.84508, 233.82309, 233.79951, 233.77438, 233.74776, 233.73389, 233.70505, 233.67479, 233.64311, 233.61003, 233.57556, 233.53972, 233.50253, 233.46399, 233.42413, 233.383, 233.34067, 233.29721, 233.25272, 233.2073, 233.16113, 233.11435, 233.06712, 233.01958, 232.97186, 232.92409, 232.8764, 232.82896, 232.78198, 232.73569, 232.69029, 232.64604, 232.6032, 232.56206, 232.52287, 232.4858, 232.46803, 232.43408, 232.4022, 232.37236, 232.34439, 232.3181, 232.29329, 232.26976, 232.24728, 232.22348, 232.20241, 232.18164, 232.16098, 232.14024, 232.11923, 232.0978, 232.07588, 232.05347, 232.0305, 232.00699, 231.99504, 231.97081, 231.94621, 231.92131, 231.89615, 231.87077, 231.8452, 231.81947, 231.79358, 231.76746, 231.74107, 231.71437, 231.68733, 231.65996, 231.63222, 231.60413, 231.57567, 231.54689, 231.51778, 231.48839, 231.45874, 231.44383, 231.41393, 231.38394, 231.35391, 231.3239, 231.29395, 231.26408, 231.23436, 231.2048, 231.17546, 231.16087, 231.13191, 231.10324, 231.07487, 231.04686, 231.0192, 230.99197, 230.96527, 230.93921, 230.91388, 230.88934, 230.86563, 230.85408, -999.0, 230.81001, 230.78911, 230.76878, 230.74887, 230.72926, 230.70985, 230.69055, 230.67131, 230.65204, 230.63272, 230.61328, 230.59373, 230.574, 230.55412, 230.53404, 230.51375, 230.49327, 230.47261, 230.46222, 230.44138, 230.42046, 230.39944, 230.37831, 230.35701, 230.33546, 230.31357, 230.2911, 230.26784, -999.0, 230.21822, 230.20514, 230.17819, 230.15025, 230.12134, 230.09163, 230.06128, 230.03046, 229.9993, 229.96785, 229.93613, 229.9041, 229.87181, 229.83928, -999.0, -999.0, -999.0, -999.0, 229.67387, 229.6403, 229.60657, 229.58624, 229.55225, 229.51811, 229.48386, 229.4495, 229.41502, 229.3805, 229.34589, 229.31117, 229.27623, 229.25865, 229.2232, 229.18729, 229.15082, 229.1137, 229.07579, 229.03706, 228.99751, 228.95718, 228.91612, 228.87434, 228.8319, 228.7888, 228.74507, 228.70078, -999.0, -999.0, -999.0, -999.0, -999.0, 228.42766, 228.40474, 228.35902, 228.31358, -999.0, -999.0, -999.0, 228.13791, 228.09636, -999.0, -999.0, 227.9803, 227.945, 227.91165, 227.88036, 227.85144, 227.82535, 227.80257, 227.78354, -999.0, 227.75597, 227.74635, 227.73877, 227.73277, 227.72795, 227.72395, 227.72038, 227.717, 227.71371, 227.71043, 227.70709, 227.70361, 227.70006, 227.69644, 227.69463, 227.69096, 227.68729, 227.6836, 227.6799}
theta =
  {310.70667, -999.0, -999.0, -999.0, -999.0, -999.0, 310.83856, 310.84335, 310.8477, 310.85147, 310.85468, 310.85736, 310.85947, 310.86105, 310.86212, 310.8627, 310.86282, 310.86258, 310.8621, 310.86154, 310.8611, 310.86096, 310.86124, 310.8621, 310.86365, 310.86606, 310.8694, 310.87363, 310.87885, 310.88504, 310.89212, 310.8999, 310.9082, 310.91684, 310.92572, 310.93463, 310.9434, 310.9519, 310.96005, 310.96783, 310.9752, 310.9821, 310.9886, 310.9947, 311.00046, 311.00598, 311.01132, 311.0166, 311.02197, 311.02756, 311.0335, 311.03995, 311.04712, 311.0551, 311.06433, 311.07504, 311.08765, 311.10245, 311.11984, 311.14017, 311.16632, 311.19394, 311.22543, 311.2611, 311.30115, 311.34576, 311.39508, 311.4491, 311.50787, 311.57138, 311.63934, 311.7114, 311.7871, 311.86606, 311.94733, 312.02988, 312.1127, 312.1949, 312.2759, 312.35535, 312.43274, 312.50775, 312.58014, 312.64984, 312.71667, 312.78043, 312.84036, 312.89575, 312.94574, 312.9897, 313.0275, 313.05923, -999.0, -999.0, -999.0, -999.0, -999.0, 313.14044, 313.14203, 313.1419, 313.1407, 313.13885, 313.1369, 313.13528, 313.1344, 313.13464, 313.13608, 313.13867, 313.14243, 313.14728, 313.15305, 313.1595, 313.16635, 313.1734, 313.18057, 313.18774, 313.19492, 313.2019, 313.20862, 313.21478, 313.22025, 313.22482, 313.22855, 313.2314, 313.23358, 313.2351, 313.2362, 313.2371, 313.23804, 313.2393, 313.24094, 313.24307, 313.24576, 313.2491, 313.25305, 313.25754, 313.26254, 313.26797, 313.2737, 313.27954, 313.28528, 313.2908, 313.29593, 313.3006, 313.30466, 313.308, 313.31073, 313.3128, 313.31433, 313.31537, 313.31604, 313.31656, 313.31702, 313.3176, 313.3183, 313.3192, 313.32028, 313.32156, 313.323, 313.3247, 313.32632, 313.32797, 313.3296, 313.33112, 313.3325, 313.3337, 313.33472, 313.3356, 313.33633, 313.33694, 313.33746, 313.33792, 313.3383, 313.3386, 313.3389, 313.3393, 313.33978, 313.34042, 313.34128, 313.34232, 313.34357, 313.345, 313.34662, 313.34827, 313.34985, 313.35135, 313.35266, 313.35373, 313.35452, 313.35492, 313.35495, 313.3546, 313.35385, 313.35266, 313.35107, 313.3491, 313.34674, 313.344, 313.34113, 313.33832, 313.33585, 313.3339, 313.33258, 313.332, 313.33228, 313.33344, 313.33557, 313.33884, 313.34326, 313.3489, 313.35568, 313.36337, 313.37177, 313.3807, 313.38998, 313.39944, 313.40894, 313.41833, 313.42764, 313.43692, 313.44623, 313.45566, 313.4654, 313.47565, 313.48666, 313.49863, 313.5116, 313.52557, 313.5406, 313.55664, 313.57358, 313.5912, 313.60922, 313.62753, 313.6459, 313.66415, 313.6821, 313.69955, 313.71637, 313.73245, 313.74762, 313.7618, 313.77487, 313.7868, 313.79752, 313.80692, 313.81497, 313.82162, 313.82684, 313.83057, 313.83286, 313.83386, 313.83365, 313.83234, 313.83008, 313.8271, 313.82352, 313.81958, 313.81537, 313.8111, 313.80685, 313.8028, 313.79898, 313.79523, 313.79224, 313.78976, 313.78778, 313.78625, 313.78513, 313.7844, 313.78384, 313.7834, 313.78284, 313.782, 313.78076, 313.779, 313.7765, 313.77316, 313.76898, 313.764, 313.7582, 313.75162, 313.74426, 313.73618, 313.7274, 313.71786, 313.70764, 313.69662, 313.68472, 313.6719, 313.65787, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 313.4468, 313.44678, 313.44577, 313.44385, 313.44095, 313.43692, 313.43158, 313.42404, 313.41553, 313.40546, 313.39374, 313.38037, 313.36563, 313.34988, 313.33353, 313.31686, 313.30023, 313.28397, 313.26834, 313.25366, 313.24, 313.22748, 313.2161, 313.206, 313.1973, 313.19022, 313.18497, 313.18167, 313.18027, 313.1806, 313.18246, 313.18573, 313.18994, 313.1947, 313.19952, 313.204, 313.2077, 313.21033, 313.21146, 313.21075, 313.2082, 313.20374, 313.19742, 313.1893, 313.1797, 313.16895, 313.1574, 313.14554, 313.13382, 313.1228, 313.11304, 313.105, 313.09906, 313.0953, 313.09396, 313.09515, 313.09897, 313.10535, 313.11432, 313.12582, 313.1396, 313.1552, 313.1724, 313.1907, 313.20975, 313.22913, 313.24835, 313.2671, 313.285, 313.3019, 313.31757, 313.3318, 313.3444, 313.3553, 313.3643, 313.37134, 313.37628, 313.37906, 313.37967, 313.37796, 313.37393, 313.36752, 313.35867, 313.34735, 313.33356, 313.31738, 313.29883, 313.27798, 313.2549, 313.2298, 313.2028, 313.174, 313.14377, 313.11234, 313.08005, 313.0472, 313.0144, 312.9822, 312.9513, 312.9195, 312.89304, 312.86932, 312.84875, 312.83163, 312.8179, 312.80743, 312.80002, 312.7955, 312.7936, 312.79398, 312.79636, 312.8004, 312.80588, 312.81253, 312.82013, 312.82843, 312.83728, 312.8465, 312.856, 312.8656, 312.87524, 312.88486, 312.8944, 312.90387, 312.91318, 312.92233, 312.93134, 312.94016, 312.94882, 312.95724, 312.9654, 312.97324, 312.98074, 312.9879, 312.99466, 313.001, 313.0069, 313.0123, 313.0172, 313.02158, 313.02536, 313.0286, 313.03122, 313.03323, 313.03464, 313.03546, 313.0357, 313.0354, 313.03458, 313.03326, 313.03152, 313.02936, 313.02682, 313.02396, 313.0208, 313.01746, 313.0139, 313.01013, 313.00616, 313.00208, 312.99783, 312.99344, 312.98898, 312.98444, 312.97992, 312.97556, 312.97147, 312.9678, 312.96472, 312.96234, 312.96088, 312.96048, 312.9612, 312.96323, 312.9666, 312.97144, 312.9779, 312.98618, 312.99646, 313.00894, 313.02386, 313.0414, 313.06183, 313.08536, 313.11206, 313.14215, 313.17566, 313.21274, 313.2534, 313.29758, 313.34528, 313.39645, 313.45102, 313.50876, 313.5695, 313.6331, 313.69907, 313.76688, 313.83603, 313.9059, 313.97598, 314.04565, 314.11435, 314.18146, 314.2466, 314.30942, 314.36954, 314.42664, 314.48065, 314.53152, 314.57928, 314.62827, 314.6696, 314.70804, 314.74365, 314.77658, 314.80685, 314.8344, 314.8593, 314.88153, 314.9009, 314.9174, 314.93082, -999.0, -999.0, -999.0, 314.9539, 314.95273, 314.94916, 314.9435, 314.93607, 314.92706, 314.9168, 314.90555, 314.8935, 314.88092, 314.86807, 314.85516, 314.8424, 314.83005, 314.81818, 314.8069, 314.7963, 314.7865, 314.77747, 314.76926, 314.76187, 314.7553, 314.7495, 314.74448, 314.74014, 314.73645, 314.7334, 314.73093, 314.729, 314.7276, 314.7267, 314.72632, 314.72644, 314.72705, 314.72815, 314.72974, 314.73184, 314.73447, 314.73758, 314.74112, 314.74506, 314.74933, 314.7538, 314.7584, 314.7629, 314.76724, 314.77133, 314.77512, 314.7785, 314.7815, 314.78406, 314.78616, 314.7878, 314.789, 314.78973, 314.79, 314.78986, 314.78925, 314.78815, 314.78644, 314.78406, 314.7809, 314.77695, 314.77206, 314.76627, 314.75943, 314.7516, 314.74274, 314.73288, 314.7221, 314.71045, 314.69806, 314.68503, 314.6715, 314.6575, 314.6431, 314.62823, 314.61145, 314.59583, 314.5799, 314.56375, 314.5474, 314.53098, 314.51453, 314.49817, 314.48196, 314.46603, 314.4506, 314.43573, 314.4216, 314.40836, 314.396, 314.38464, 314.37433, 314.36493, 314.35626, 314.34814, 314.34033, 314.33255, 314.32446, 314.31573, 314.30603, 314.29547, 314.28424, 314.27264, 314.2609, 314.24927, 314.23807, 314.22763, 314.2182, 314.2098, 314.2025, 314.1962, 314.19086, 314.18616, 314.18173, 314.17715, 314.17206, 314.1662, 314.1595, 314.15182, 314.14304, 314.13315, 314.12216, 314.11005, 314.09683, 314.08273, 314.06808, 314.05316, 314.03824, 314.02368, 314.00977, 313.9968, 313.98508, 313.9749, 313.96658, 313.96036, 313.95654, 313.9554, 313.9572, 313.96222, 313.97067, 313.9827, 313.9983, 314.0175, 314.04028, 314.06613, 314.09418, 314.12357, 314.15353, 314.1834, 314.2127, 314.2409, 314.2676, 314.29282, 314.3169, 314.34024, 314.36325, 314.38623, 314.40964, 314.43387, 314.45926, 314.48584, 314.51343, 314.5419, 314.57108, 314.6006, 314.6301, 314.6592, 314.68756, 314.7151, 314.7418, 314.76776, 314.79306, 314.81772, 314.84177, 314.8653, 314.8883, 314.9109, 314.93527, 314.95718, 314.97885, 315.00024, 315.0213, 315.04187, 315.0619, 315.08127, 315.09988, 315.11765, 315.1345, 315.15036, 315.16528, 315.17923, 315.1922, 315.2042, 315.21518, 315.22522, 315.23425, 315.24237, 315.24966, 315.25623, 315.26218, 315.26764, 315.27277, 315.27777, 315.2828, 315.28806, 315.29364, 315.2997, 315.30646, 315.31396, 315.32227, 315.33145, 315.3416, 315.3527, 315.36465, 315.37747, 315.3911, 315.40543, 315.42038, 315.43576, 315.4515, 315.46747, 315.48346, 315.49933, 315.51486, 315.52994, 315.54443, 315.55814, 315.57098, 315.58292, 315.58856, 315.59927, 315.60925, 315.6186, 315.62738, 315.63574, 315.64383, 315.65176, 315.6596, 315.66745, 315.67545, 315.6836, 315.69196, 315.70056, 315.7094, 315.7185, 315.72775, 315.73703, 315.74625, 315.7553, 315.76407, 315.77252, 315.78052, 315.78802, 315.7949, 315.80106, 315.80646, 315.811, 315.81482, 315.81796, 315.8206, 315.82278, 315.82468, 315.8264, 315.82803, 315.82977, 315.8318, 315.8342, 315.83725, 315.84106, 315.84583, 315.85175, 315.85895, 315.8676, 315.8778, 315.88962, 315.90308, 315.91827, 315.93515, 315.95358, 315.9756, 315.99713, 316.02002, 316.04425, 316.0697, 316.09637, 316.1242, 316.15323, 316.18335, 316.21463, 316.24707, 316.28073, 316.31564, 316.35184, 316.38913, 316.4274, 316.4665, 316.50616, 316.54602, 316.5856, 316.6245, 316.66232, 316.69864, 316.73315, 316.7655, 316.7954, 316.82278, 316.8476, 316.86975, 316.88928, 316.90643, 316.92136, 316.9343, 316.94553, 316.95535, 316.96408, 316.97208, 316.97958, 316.98697, 316.99445, 317.0023, 317.01077, 317.01996, 317.02994, 317.04077, 317.05252, 317.0651, 317.07846, 317.0925, 317.10712, 317.12198, 317.13672, 317.15103, 317.16455, 317.17703, 317.18808, 317.19748, 317.20502, 317.21072, 317.21472, 317.2171, 317.218, 317.21762, 317.21628, 317.21414, 317.21143, 317.2083, 317.20486, 317.20123, 317.19754, 317.19385, 317.19028, 317.18692, 317.1838, 317.18097, 317.17847, 317.17627, 317.17438, 317.17282, 317.17154, 317.17053, 317.1698, 317.16934, 317.1692, 317.16937, 317.16986, 317.1707, 317.17184, 317.17334, 317.17514, 317.17725, 317.17957, 317.182, 317.1846, 317.18726, 317.19, 317.19287, 317.19577, 317.19882, 317.20197, 317.20526, 317.20868, 317.21252, 317.21597, 317.2193, 317.2224, 317.22522, 317.22766, 317.2296, 317.23105, 317.23196, 317.2323, 317.2321, 317.23132, 317.22998, 317.22803, 317.2255, 317.22238, 317.2187, 317.21457, 317.21008, 317.2053, 317.20044, 317.19568, 317.19128, 317.18747, 317.1846, 317.18295, 317.18295, 317.18488, 317.18896, 317.19556, 317.2048, 317.217, 317.23233, 317.25095, 317.27298, 317.29868, 317.32803, 317.36124, 317.39835, 317.43942, 317.48447, 317.50848, 317.55942, 317.61423, 317.67276, 317.73474, 317.7999, 317.86795, 317.9386, 318.0114, 318.08606, 318.1621, 318.2392, 318.31686, 318.39468, 318.47226, 318.549, 318.6244, 318.6978, 318.7687, 318.83655, 318.90085, 318.9611, 319.01678, 319.06775, 319.11395, 319.15536, 319.19196, 319.2239, 319.2515, 319.275, 319.2947, 319.3109, 319.32404, 319.33435, 319.34225, 319.34805, 319.35214, 319.3548, 319.3564, 319.35736, 319.35797, 319.3587, 319.3599, 319.3619, 319.36502, 319.3695, 319.37564, 319.38364, 319.3936, 319.40555, 319.41965, 319.43585, 319.45413, 319.47433, 319.49643, 319.5203, 319.5457, 319.57242, 319.60034, 319.6293, 319.65912, 319.68973, 319.72095, 319.75266, 319.78467, 319.81677, 319.84885, 319.88058, 319.9118, 319.94223, 319.9716, 319.99973, 320.02914, 320.05444, 320.07828, 320.10062, 320.12158, 320.14117, 320.15952, 320.1766, 320.19263, 320.20758, 320.22162, 320.23486, 320.2474, 320.25937, 320.27094, 320.28217, 320.29315, 320.30402, 320.31482, 320.32562, 320.33646, 320.3419, 320.3528, 320.36377, 320.37476, 320.38574, 320.39673, 320.40762, 320.41837, 320.4289, 320.43915, 320.44904, 320.4586, 320.46774, 320.47647, 320.4848, 320.49274, 320.50034, 320.50763, 320.51465, 320.5214, 320.52798, 320.53442, 320.54074, 320.547, 320.55322, 320.55945, 320.56573, 320.57208, 320.57846, 320.5849, 320.59137, 320.5978, 320.6042, 320.6104, 320.61642, 320.62228, 320.62793, 320.63342, 320.63876, 320.64398, 320.64908, 320.6541, 320.65912, 320.66406, 320.66895, 320.67377, 320.67847, 320.68314, 320.68777, 320.69244, 320.69714, 320.70197, 320.70694, 320.71216, 320.71762, 320.72342, 320.72958, 320.7361, 320.7431, 320.7505, 320.75824, 320.76636, 320.77478, 320.78348, 320.79248, 320.80173, 320.81125, 320.82104, 320.83127, 320.84198, 320.85327, 320.86523, 320.878, 320.89166, 320.9063, 320.92197, 320.93854, 320.956, 320.97427, 320.99323, 321.0126, 321.03223, 321.04404, 321.06363, 321.083, 321.102, 321.12042, 321.13818, 321.15518, 321.1713, 321.1865, 321.20065, 321.21368, 321.22552, 321.23608, 321.2454, 321.25357, 321.26068, 321.2668, 321.2722, 321.277, 321.28152, 321.28595, 321.29053, 321.29535, 321.30066, 321.30658, 321.3132, 321.3206, 321.32874, 321.33774, 321.34756, 321.3583, 321.36996, 321.38263, 321.39633, 321.4111, 321.42697, 321.444, 321.46216, 321.48145, 321.50177, 321.5231, 321.5454, 321.56866, 321.59283, 321.6179, 321.6439, 321.6708, 321.6987, 321.72763, 321.75757, 321.78842, 321.8201, 321.85254, 321.88562, 321.9192, 321.9531, 321.98718, 322.02115, 322.0547, 322.08743, 322.12784, 322.15814, 322.1869, 322.2139, 322.23907, 322.26242, 322.28406, 322.30417, 322.32294, 322.34055, 322.3571, 322.37277, 322.38773, 322.40213, 322.41614, 322.42993, 322.44363, 322.4575, 322.4717, 322.48654, 322.5022, 322.51892, 322.52774, 322.54645, 322.56668, 322.58868, 322.61243, 322.63788, 322.66498, 322.69373, 322.72385, 322.75513, 322.79056, 322.82346, 322.85666, 322.88992, 322.92294, 322.95538, 322.98715, 323.01804, 323.04785, 323.07648, 323.10382, 323.12985, 323.15445, 323.17764, 323.19937, 323.21973, 323.2387, 323.25635, 323.27267, 323.2878, 323.30173, 323.3145, 323.3261, 323.3365, 323.3456, 323.35342, 323.35977, 323.36453, 323.36752, 323.3686, 323.36755, 323.36426, 323.35852, 323.3502, 323.3394, 323.32623, 323.31085, 323.2935, 323.2746, 323.25467, 323.23425, 323.21387, 323.194, 323.17514, 323.15784, 323.14255, 323.12958, 323.11932, 323.1121, 323.10812, 323.10748, 323.10837, 323.1126, 323.12006, 323.13055, 323.1438, 323.15955, 323.17752, 323.19745, 323.21902, 323.242, 323.2661, 323.29126, 323.31744, 323.34464, 323.3729, 323.40234, 323.43314, 323.46545, 323.4995, 323.53555, 323.5738, 323.6145, 323.658, 323.7044, 323.7539, 323.80655, 323.8625, 323.9216, 323.98367, 324.0484, 324.11554, 324.18472, 324.25558, 324.32773, 324.40076, 324.47424, 324.54785, 324.62112, 324.6937, 324.76517, 324.83524, 324.90353, 324.93695, 325.00204, 325.06482, 325.1252, 325.1832, 325.23877, 325.292, 325.343, 325.39188, 325.4388, 325.4883, 325.53143, 325.5729, 325.6128, 325.65115, 325.688, 325.72336, 325.7573, 325.78976, 325.82083, 325.85043, 325.8786, 325.90536, 325.93066, 325.9545, 325.9769, 325.99786, 326.01746, 326.03568, 326.05252, 326.0681, 326.0824, 326.0955, 326.10733, 326.118, 326.12753, 326.13596, 326.14325, 326.1495, 326.15485, 326.15936, 326.16312, 326.1662, 326.1687, 326.17075, 326.17242, 326.17392, 326.17538, 326.17706, 326.17908, 326.1817, 326.18524, 326.18994, 326.196, 326.20358, 326.2128, 326.22375, 326.23648, 326.25095, 326.2671, 326.28485, 326.30408, 326.32468, 326.3464, 326.36914, 326.3927, 326.4169, 326.44156, 326.46652, 326.49158, 326.5167, 326.5418, 326.5668, 326.5916, 326.61627, 326.64072, 326.6649, 326.68884, 326.71243, 326.73563, 326.75836, 326.78055, 326.80215, 326.82318, 326.84366, 326.86353, 326.88287, 326.9018, 326.92038, 326.93872, 326.95685, 326.97485, 326.9927, 327.01053, 327.0283, 327.04602, 327.06372, 327.08148, 327.09927, 327.11713, 327.13507, 327.15314, 327.16223, 327.18042, 327.19867, 327.21692, 327.23514, 327.25323, 327.27118, 327.2889, 327.30634, 327.3235, 327.34198, 327.3584, 327.37445, 327.39014, 327.40543, 327.42035, 327.4349, 327.44916, 327.46307, 327.47678, 327.49023, 327.50357, 327.51685, 327.5301, 327.5434, 327.55664, 327.5699, 327.58304, 327.59607, 327.60898, 327.6217, 327.63422, 327.64645, 327.65842, 327.66998, 327.68118, 327.69193, 327.70212, 327.71173, 327.7207, 327.7289, 327.73636, 327.743, 327.74875, 327.75363, 327.75763, 327.76077, 327.76306, 327.76453, 327.76517, 327.76505, 327.76413, 327.76248, 327.76013, 327.7571, 327.7535, 327.74936, 327.74475, 327.73975, 327.73447, 327.729, 327.7235, 327.71817, 327.71313, 327.70865, 327.705, 327.7025, 327.70154, 327.70276, 327.70728, 327.71625, 327.73083, 327.75125, 327.77667, 327.8062, 327.83896, 327.87405, 327.9106, 327.94772, 327.98456, 328.0205, 328.05542, 328.07245, 328.10547, 328.13702, 328.1672, 328.1961, 328.22385, 328.25052, 328.27634, 328.30142, 328.32605, 328.3503, 328.37448, 328.3987, 328.42322, 328.44818, 328.47366, 328.49973, 328.52643, 328.55377, 328.58173, 328.6101, 328.6389, 328.66794, 328.69708, 328.7262, 328.75513, 328.7837, 328.8117, 328.83887, 328.86493, 328.88965, 328.91296, 328.93484, 328.9553, 328.97427, 328.99197, 329.0085, 329.02408, 329.03882, 329.05286, 329.0663, 329.08054, 329.09305, 329.10526, 329.11722, 329.1291, 329.14093, 329.1528, 329.16476, 329.17685, 329.1891, 329.2015, 329.2141, 329.2269, 329.2398, 329.2529, 329.2661, 329.27945, 329.29294, 329.30652, 329.3202, 329.33398, 329.34787, 329.36185, 329.37592, 329.3901, 329.40442, 329.4188, 329.43323, 329.4477, 329.46213, 329.47656, 329.49112, 329.50577, 329.5206, 329.53564, 329.5509, 329.5664, 329.58218, 329.59827, 329.61462, 329.6313, 329.6483, 329.66562, 329.6833, 329.7013, 329.71964, 329.73828, 329.7572, 329.77634, 329.79572, 329.81522, 329.83484, 329.8545, 329.87415, 329.89377, 329.91327, 329.93268, 329.9519, 329.97095, 329.9898, 330.0084, 330.0268, 330.04498, 330.06308, 330.08112, 330.0992, 330.11743, 330.13602, 330.15503, 330.17465, 330.195, 330.21622, 330.23843, 330.26175, 330.28635, 330.31226, 330.3397, 330.36868, 330.3994, 330.43195, 330.46634, 330.50275, 330.54105, 330.58115, 330.62292, 330.66626, 330.71085, 330.75644, 330.80267, 330.84927, 330.8959, 330.94226, 330.98798, 331.03278, 331.0762, 331.1179, 331.15738, 331.19427, 331.22836, 331.25943, 331.2873, 331.31183, 331.33496, 331.3527, 331.36734, 331.3791, 331.38812, 331.3947, 331.3991, 331.40155, 331.40228, 331.40152, 331.39957, 331.39667, 331.39307, 331.38904, 331.38486, 331.38077, 331.377, 331.37375, 331.37112, 331.36932, 331.36844, 331.3685, 331.36957, 331.37167, 331.3747, 331.3785, 331.38287, 331.38763, 331.3926, 331.39755, 331.40222, 331.4064, 331.41006, 331.41327, 331.41595, 331.4182, 331.42004, 331.42154, 331.42273, 331.42368, 331.42438, 331.42487, 331.42514, 331.4252, 331.4251, 331.42496, 331.42474, 331.42456, 331.42438, 331.42413, 331.4238, 331.42337, 331.42282, 331.4222, 331.42163, 331.42114, 331.42078, 331.4207, 331.4209, 331.42157, 331.4227, 331.42432, 331.4265, 331.42932, 331.43268, 331.43665, 331.44116, 331.44623, 331.45178, 331.45776, 331.46408, 331.47064, 331.47742, 331.48087, 331.48776, 331.4947, 331.50156, 331.50833, 331.51492, 331.52133, 331.52744, 331.53333, 331.5389, 331.54163, 331.5468, 331.55185, 331.55685, 331.562, 331.56744, 331.5732, 331.57944, 331.58615, 331.5934, 331.60196, 331.6102, 331.61877, 331.62762, 331.6367, 331.64587, 331.65518, 331.66452, 331.67392, 331.6834, 331.69302, 331.70276, 331.71268, 331.72284, 331.73334, 331.74417, 331.7554, 331.76697, 331.77893, 331.79123, 331.79745, 331.80994, 331.82233, 331.83444, 331.84598, 331.8566, 331.8659, 331.8736, 331.8792, 331.88242, 331.88278, 331.88177, 331.87717, 331.869, 331.85715, 331.84155, 331.82217, 331.79916, 331.77274, 331.74313, 331.71066, 331.67575, 331.65756, 331.62003, 331.58145, 331.54236, 331.50342, 331.46518, 331.42825, 331.39328, 331.3608, 331.33148, 331.30582, 331.28442, 331.26785, 331.2566, 331.25122, 331.25253, 331.26166, 331.27985, 331.30832, 331.3473, 331.39532, 331.4509, 331.51242, 331.57812, 331.646, 331.7139, 331.77972, 331.84195, 331.89993, 331.95312, 332.001, 332.04324, 332.07993, 332.1111, 332.137, 332.15775, 332.17383, 332.18567, 332.1938, 332.19864, 332.20068, 332.20044, 332.1996, 332.19678, 332.19284, 332.18814, 332.18317, 332.17825, 332.1737, 332.1697, 332.16644, 332.16412, 332.1634, 332.16278, 332.16354, 332.1658, 332.16965, 332.17505, 332.18204, 332.19052, 332.20053, 332.21198, 332.22482, 332.23178, 332.24667, 332.26282, 332.28015, 332.29852, 332.31787, 332.3381, 332.35913, 332.38086, 332.39197, 332.41467, 332.42856, 332.4522, 332.4764, 332.5012, 332.52643, 332.552, 332.57776, 332.60358, 332.62927, 332.65457, 332.67923, 332.70306, 332.72604, 332.74823, 332.76968, 332.7905, 332.81067, 332.83035, 332.84958, 332.86844, 332.88705, 332.9056, 332.92422, 332.9431, 332.9624, 332.98224, 333.0028, 333.02423, 333.04663, 333.0702, 333.09497, 333.10785, 333.1347, 333.16293, 333.19257, 333.22363, 333.2561, 333.28992, 333.325, 333.3613, 333.39865, 333.43677, 333.47537, 333.51416, 333.55273, 333.59058, 333.62708, 333.66168, 333.69388, 333.72318, 333.74905, 333.77112, 333.78906, 333.80286, 333.81262, 333.8184, 333.82047, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 335.25806, 335.28714, 335.3103, 335.32684, 335.33597, 335.33698, 335.3298, 335.3159, 335.29684, 335.27417, 335.24927, 335.223, 335.19617, 335.16956, 335.1439, 335.11957, 335.09695, 335.07645, 335.0583, 335.04254, 335.02924, 335.01834, 335.00992, 335.00378, 334.99985, 334.998, 334.99805, 334.99988, 335.0032, 335.0079, 335.0137, 335.02036, 335.0276, 335.0351, 335.04263, 335.04996, 335.05692, 335.06323, 335.0688, 335.07333, 335.07672, 335.07874, 335.07916, 335.07895, 335.07733, 335.0744, 335.0702, 335.06485, 335.05853, 335.05145, 335.0437, 335.0355, 335.02686, 335.01794, 335.0088, 334.9995, 334.99014, 334.9807, 334.97125, 334.96176, 334.95215, 334.94238, 334.93237, 334.9273, 334.91708, 334.90683, 334.89667, 334.88672, 334.87723, 334.86835, 334.8603, 334.85324, 334.8473, 334.84256, 334.8391, 334.83704, 334.83627, 334.83676, 334.83847, 334.8413, 334.84515, 334.8498, 334.85507, 334.86087, 334.8671, 334.87372, 334.88068, 334.88794, 334.89557, 334.9035, 334.91187, 334.9206, 334.92975, 334.94037, 334.9505, 334.96112, 334.97214, 334.9835, 334.99506, 335.0068, 335.0186, 335.03036, 335.04202, 335.0535, 335.06482, 335.076, 335.08707, 335.09805, 335.10892, 335.11966, 335.13025, 335.14072, 335.15103, 335.1612, 335.17123, 335.17624, 335.1861, 335.1958, 335.20538, 335.21475, 335.2239, 335.23282, 335.24142, 335.24966, 335.2575, 335.26495, 335.27197, 335.27856, 335.2847, 335.29047, 335.29587, 335.301, 335.30585, 335.31052, 335.31503, 335.31943, 335.32373, 335.32806, 335.3324, 335.33682, 335.34146, 335.34647, 335.352, 335.35822, 335.3652, 335.37308, 335.38184, 335.38657, 335.39676, 335.4078, 335.41962, 335.43213, 335.44513, 335.4585, 335.472, 335.48538, 335.49197, 335.50473, 335.5167, 335.52756, 335.537, 335.5448, 335.5509, 335.5552, 335.55765, 335.5582, 335.55692, 335.5556, 335.5517, 335.54605, 335.53873, 335.52966, 335.51886, 335.50638, 335.49265, 335.47797, 335.4628, 335.44757, 335.4401, 335.4258, 335.41296, 335.4021, 335.39395, 335.38934, 335.38904, 335.3939, 335.40424, 335.4221, 335.44427, 335.47217, 335.50464, 335.54016, 335.577, 335.61362, 335.64917, 335.6832, 335.71533, 335.74515, 335.7725, 335.78525, 335.8089, 335.83008, 335.84888, 335.8656, 335.88052, 335.89395, 335.90616, 335.91733, 335.92758, 335.9371, 335.94162, 335.95016, 335.95798, 335.965, 335.97116, 335.97644, 335.98077, 335.9842, 335.9866, 335.98804, 335.98856, 335.98846, 335.9876, 335.98584, 335.98322, 335.9797, 335.9753, 335.97006, 335.96396, 335.957, 335.94922, 335.945, 335.93594, 335.92587, 335.9147, 335.90234, 335.88885, 335.87445, 335.85934, 335.84372, 335.8279, 335.81232, 335.7973, 335.7833, 335.7711, 335.76172, 335.75623, 335.7556, 335.7603, 335.7703, 335.7855, 335.80582, 335.81775, 335.8443, 335.8735, 335.90424, 335.9355, 335.96692, 335.9983, 336.0294, 336.05997, 336.09003, 336.1195, 336.14838, 336.17664, 336.20444, 336.23187, 336.2591, 336.2863, 336.31342, 336.34055, 336.3677, 336.39484, 336.4219, 336.44876, 336.47522, 336.50122, 336.52658, 336.5511, 336.57462, 336.59692, 336.61783, 336.6371, 336.646, 336.66232, 336.67654, 336.68866, 336.6987, 336.70663, 336.7126, 336.71667, 336.71915, 336.72012, 336.7201, 336.71918, 336.71722, 336.71445, 336.711, 336.7071, 336.7028, 336.6983, 336.69373, 336.6892, 336.68448, 336.68054, 336.6771, 336.67435, 336.67242, 336.67157, 336.67188, 336.67346, 336.67645, 336.68088, 336.68686, 336.69043, 336.69873, 336.70856, 336.7199, 336.73276, 336.74704, 336.76263, 336.7795, 336.79755, 336.81665, 336.83676, 336.84717, 336.86862, 336.89102, 336.9145, 336.9391, 336.96497, 336.99228, 337.02118, 337.0519, 337.08463, 337.11935, 337.13745, 337.17526, 337.21515, 337.257, 337.3005, 337.3454, 337.39142, 337.43817, 337.48517, 337.53198, 337.57812, 337.60083, 337.64536, 337.68854, 337.7301, 337.7699, 337.80792, 337.8442, 337.87878, 337.91174, 337.94305, 337.97275, 337.98703, 338.0144, 338.04016, 338.0642, 338.0865, 338.1069, 338.1253, 338.14157, 338.15558, 338.16718, 338.17633, 338.18298, 338.18716, 338.18884, 338.1881, 338.1852, 338.18027, 338.17352, 338.16522, 338.1557, 338.14523, 338.13412, 338.1228, 338.1117, 338.10126, 338.09192, 338.08417, 338.07843, 338.07513, 338.07468, 338.0773, 338.07977, 338.087, 338.09735, 338.1107, 338.12677, 338.1453, 338.16586, 338.18817, 338.21185, 338.23904, 338.2644, 338.29007, 338.3157, 338.3411, 338.366, 338.39017, 338.41357, 338.4362, 338.45804, 338.47903, 338.48923, 338.50903, 338.52808, 338.54633, 338.56384, 338.5806, 338.59665, 338.612, 338.62665, 338.64056, 338.65372, 338.66608, 338.6776, 338.68826, 338.69788, 338.70645, 338.71396, 338.72055, 338.7263, 338.73132, 338.73575, 338.7378, 338.74164, 338.7453, 338.74893, 338.7527, 338.75674, 338.76123, 338.7663, 338.772, 338.77844, 338.78195, 338.78955, 338.798, 338.8073, 338.81747, 338.82852, 338.84048, 338.85342, 338.8673, 338.88226, 338.89813, 338.9149, 338.92352, 338.94128, 338.95956, 338.9782, 338.99707, 339.016, 339.03482, 339.05347, 339.07184, 339.08994, 339.1076, 339.12488, 339.14166, 339.15793, 339.1737, 339.18903, 339.204, 339.21875, 339.23334, 339.24786, 339.25516, 339.26987, 339.2848, 339.30002, 339.31552, 339.3313, 339.34735, 339.36353, 339.37967, 339.3956, 339.41107, 339.42606, 339.43338, 339.44766, 339.46158, 339.4751, 339.4883, 339.50128, 339.51404, 339.52667, 339.5391, 339.55127, 339.5632, 339.57477, 339.58594, 339.59665, 339.6068, 339.6164, 339.62537, 339.63373, 339.6415, 339.6487, 339.65277, 339.65915, 339.66504, 339.67056, 339.67566, 339.68024, 339.68417, 339.68738, 339.68973, 339.69104, 339.69125, 339.6907, 339.68875, 339.68533, 339.68042, 339.67395, 339.66592, 339.6565, 339.64575, 339.6338, 339.6208, 339.6068, 339.592, 339.57648, 339.56033, 339.54373, 339.53616, 339.51935, 339.50262, 339.4861, 339.46997, 339.46204, 339.4466, 339.43182, 339.41782, 339.40475, 339.39276, 339.38202, 339.37262, 339.3647, 339.3583, 339.35373, 339.3512, 339.351, 339.35342, 339.359, 339.36856, 339.38284, 339.4026, -999.0, 339.4576, 339.49127, 339.5279, 339.56677, 339.60724, 339.64862, 339.69025, 339.73175, 339.77298, 339.81378, 339.854, 339.89365, 339.93283, 339.97162, 339.99088, 340.02927, 340.0675, 340.10562, 340.1437}
theta_e =
  {350.7142, -999.0, -999.0, -999.0, -999.0, -999.0, 349.31183, 349.19867, 349.0857, 348.97263, 348.86142, 348.75275, 348.64462, 348.53738, 348.43173, 348.32846, 348.2284, 348.1324, 348.0416, 347.95718, 347.88116, 347.81586, 347.76013, 347.71497, 347.68134, 347.6602, 347.6522, 347.65805, 347.67834, 347.71353, 347.76318, 347.82663, 347.90317, 347.992, 348.09164, 348.2005, 348.31702, 348.4417, 348.57123, 348.70273, 348.83417, 348.96344, 349.0884, 349.20697, 349.317, 349.4167, 349.5058, 349.58438, 349.6525, 349.71027, 349.7575, 349.79413, 349.81995, 349.83475, 349.8382, 349.82993, -999.0, 349.77664, 349.7323, 349.67764, 349.60703, 349.53424, 349.4532, 349.36334, 349.2642, 349.15744, 349.04376, 348.91962, 348.78445, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 346.32928, -999.0, -999.0, -999.0, 345.14728, 344.84464, 344.53613, 344.22772, 343.91852, 343.60297, 343.2903, 342.97495, -999.0, -999.0, -999.0, -999.0, -999.0, 341.11893, 340.8314, 340.55975, 340.29517, 340.03778, 339.79233, 339.5568, -999.0, 339.10504, 338.89526, 338.6925, 338.49628, 338.30667, 338.12952, 337.95883, 337.7939, 337.63458, -999.0, -999.0, 337.20572, 337.07587, 336.95224, 336.83643, 336.72937, 336.6281, 336.53262, 336.4428, 336.3586, 336.27988, 336.2073, 336.14154, 336.08038, 336.02362, 335.97107, 335.92264, 335.87817, 335.83762, 335.80127, 335.7696, 335.74292, 335.72165, 335.7057, 335.69495, 335.6892, 335.68854, 335.69205, 335.6988, 335.70804, 335.719, 335.73083, 335.74258, 335.7534, 335.76233, 335.7687, 335.77188, 335.77118, 335.76614, 335.75723, 335.74527, 335.731, 335.71518, 335.69843, 335.67957, 335.66257, 335.64633, 335.63132, 335.6181, 335.6072, 335.59915, 335.5942, 335.59274, 335.59497, 335.60104, 335.61038, 335.6222, 335.63568, 335.65002, 335.66443, 335.67792, 335.68967, 335.69885, 335.7051, 335.70813, 335.70764, 335.70343, 335.69528, 335.68317, 335.667, 335.64655, 335.62158, 335.59167, 335.5565, 335.51584, 335.47055, 335.4217, 335.37238, 335.32175, 335.27097, 335.22116, 335.17346, 335.12894, 335.08804, 335.05112, 335.01852, 334.9903, 334.96515, 334.94144, 334.91745, 334.89166, 334.8634, 334.83286, 334.7998, 334.7631, 334.72302, 334.68005, 334.63464, 334.58725, 334.5381, 334.4873, 334.435, 334.38138, 334.32648, 334.2728, 334.21805, 334.16232, 334.10602, 334.0496, 333.99347, 333.93814, 333.8838, 333.8307, 333.78033, 333.7328, 333.6869, 333.6427, 333.6002, 333.5593, 333.51926, 333.479, 333.43753, 333.39386, 333.34885, 333.30066, 333.2478, 333.18967, 333.12665, 333.05957, 332.9892, 332.91644, 332.84442, 332.7737, 332.70468, 332.63858, 332.5762, 332.51813, 332.46484, 332.41684, 332.37418, 332.33676, 332.30484, 332.2785, 332.25714, 332.2409, 332.22998, 332.22467, 332.22595, 332.2365, 332.25574, 332.2854, 332.32678, 332.38214, 332.45135, 332.5352, 332.63376, 332.74695, 332.87463, 333.01736, 333.17776, 333.3509, 333.5357, 333.73346, 333.945, 334.1645, 334.39188, -999.0, -999.0, 335.12042, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 334.6033, 334.47983, 334.36105, 334.2478, 334.13068, 334.03204, 333.9433, 333.86212, 333.78885, 333.72333, 333.66525, 333.6143, 333.57007, 333.53214, 333.49994, 333.47296, -999.0, -999.0, 333.4155, 333.40045, 333.38562, 333.37033, -999.0, -999.0, -999.0, -999.0, 333.27283, 333.2462, 333.2159, 333.18198, 333.14426, 333.10278, 333.05756, 333.0088, 332.95682, 332.90195, 332.84448, 332.78662, 332.72717, 332.66602, 332.60358, 332.54077, 332.47876, 332.41864, 332.36166, 332.30923, 332.26294, 332.22424, 332.19467, 332.17505, 332.16647, 332.1689, 332.18292, 332.20883, 332.2473, 332.29807, 332.36108, 332.43567, 332.52084, 332.61563, 332.719, 332.82944, 332.94516, 333.06454, 333.1875, 333.31296, 333.4384, 333.56284, 333.6854, 333.8051, 333.92105, 334.03357, 334.14227, 334.24454, 334.33975, 334.4273, 334.50665, 334.57764, 334.6403, 334.69464, 334.74078, 334.7793, 334.81143, 334.83646, 334.85495, 334.8679, 334.87646, 334.8819, 334.88525, 334.88712, 334.8878, 334.88763, 334.88702, 334.88666, 334.88736, 334.89005, -999.0, -999.0, 334.9197, 334.93878, 334.96362, 334.9941, 335.0298, 335.0703, 335.1151, 335.1629, 335.21207, 335.26105, 335.3085, 335.35397, 335.39752, 335.4391, 335.47888, 335.5171, 335.55386, 335.5896, 335.62463, 335.65942, 335.69446, 335.73013, 335.76694, 335.80496, 335.84424, 335.88477, 335.92654, 335.96933, 336.01273, 336.05643, 336.10004, 336.14264, -999.0, -999.0, 336.25354, 336.28168, 336.30417, 336.3203, 336.32953, 336.3318, 336.3273, 336.3163, 336.299, 336.27594, 336.2477, 336.2164, 336.18155, 336.14377, 336.10394, 336.06302, 336.02182, 335.98108, 335.9414, 335.90335, 335.86752, 335.83395, 335.8026, 335.7734, 335.74622, 335.72095, 335.6974, 335.67648, 335.657, 335.63867, 335.62112, 335.60413, 335.5874, 335.57095, 335.55484, 335.53918, 335.52408, 335.50974, 335.49634, 335.48422, 335.4735, 335.46402, 335.45532, 335.44708, 335.43887, 335.43, 335.41974, 335.4073, 335.39297, 335.3762, 335.35532, 335.32962, -999.0, -999.0, 335.21857, 335.16956, -999.0, -999.0, -999.0, -999.0, -999.0, 334.77304, 334.6907, -999.0, -999.0, 334.39957, 334.2927, 334.17877, -999.0, -999.0, 333.8166, -999.0, 333.57193, 333.45593, 333.3432, 333.23553, 333.1309, 333.0442, 332.96643, 332.8986, 332.84247, 332.7991, 332.76514, 332.7399, 332.7225, 332.71185, 332.7066, 332.70538, -999.0, -999.0, -999.0, 332.72025, 332.72543, 332.73016, 332.73413, 332.73694, 332.73834, 332.73834, 332.73706, 332.73456, 332.73108, 332.72748, 332.72495, 332.72467, 332.72772, 332.73517, 332.748, 332.7671, 332.79337, 332.82703, 332.86804, 332.91632, 332.9717, 333.03317, 333.09927, 333.16953, 333.2431, 333.3173, 333.3908, 333.4624, 333.5309, 333.5958, -999.0, -999.0, -999.0, 333.81195, 333.854, 333.89148, 333.92334, 333.95007, 333.97256, 333.99167, 334.0082, 334.02274, 334.03564, 334.0473, 334.05804, 334.06775, 334.07596, 334.0823, -999.0, -999.0, 334.0872, 334.08377, 334.07776, 334.06937, 334.0591, 334.0478, 334.03516, 334.02112, 334.00546, 333.98788, 333.96805, 333.94547, 333.91953, -999.0, 333.85504, 333.81604, 333.77304, 333.72647, 333.67682, 333.62476, 333.57104, 333.5164, 333.4616, 333.40826, 333.3564, 333.3059, 333.25247, 333.2061, 333.16196, 333.12018, 333.08087, 333.0437, 333.00818, 332.9738, 332.9401, 332.90698, 332.87457, 332.84293, 332.81213, 332.7824, 332.7541, 332.7274, 332.70258, 332.6795, 332.658, 332.6378, 332.61874, 332.60086, 332.5833, 332.5657, 332.54776, 332.5297, 332.5121, 332.4954, 332.48016, 332.4666, 332.45477, 332.44476, 332.43665, 332.4302, 332.42508, 332.42096, 332.4174, 332.41367, 332.40884, 332.40198, 332.3922, 332.37918, 332.36276, 332.34286, 332.3194, 332.2922, 332.26114, 332.226, 332.18677, 332.144, 332.09875, 332.052, 332.00473, 331.9577, 331.91293, 331.86996, 331.82925, 331.79132, 331.75644, 331.72504, 331.69745, 331.6744, 331.65683, 331.64563, 331.6417, 331.6458, 331.65875, 331.68127, 331.71396, 331.75616, 331.80652, 331.8636, 331.926, 331.99255, 332.0623, 332.13406, 332.20697, 332.28067, 332.3552, 332.4307, 332.50723, 332.5853, 332.66553, 332.74908, 332.83728, 332.9288, 333.02307, 333.1195, 333.21738, 333.31528, 333.4112, 333.5032, 333.58945, 333.6692, 333.74234, 333.8088, 333.86856, 333.9217, 333.96844, 334.00903, 334.04367, 334.0727, 334.0986, 334.11716, 334.13132, 334.1417, 334.14896, 334.1538, 334.15692, 334.15884, 334.16028, 334.16174, 334.16388, 334.16693, 334.17105, 334.17636, 334.18298, 334.19086, 334.19977, 334.20956, 334.22003, 334.231, 334.24216, 334.2534, 334.26443, 334.27518, 334.2855, 334.2953, 334.3045, 334.3129, 334.3202, 334.32617, 334.33054, 334.33322, 334.3341, 334.3332, 334.33038, 334.32584, 334.31976, 334.31235, 334.30383, 334.29428, 334.28378, 334.27246, 334.2603, 334.2475, 334.23514, 334.2225, 334.20953, 334.1964, 334.1833, 334.17038, 334.15784, 334.14578, 334.13998, 334.1289, 334.11856, 334.10907, 334.10037, 334.0924, 334.08514, 334.0785, 334.07233, 334.06653, 334.06097, 334.0556, 334.05063, 334.0463, 334.04288, 334.04053, 334.03934, 334.03943, 334.04086, 334.04358, 334.0472, 334.05136, 334.0557, 334.06006, 334.06403, 334.0674, 334.07007, 334.07187, 334.0727, 334.0725, 334.07117, 334.06857, 334.0645, 334.05875, -999.0, -999.0, 334.02997, 334.017, 334.00284, 333.9878, 333.97247, 333.95746, 333.94333, 333.93076, 333.92023, 333.9124, 333.90784, 333.90695, 333.90985, 333.9166, 333.9285, 333.9433, 333.96164, 333.98322, 334.00778, 334.03494, 334.0642, 334.09543, 334.12775, 334.1607, 334.19394, 334.22714, 334.25998, 334.29214, -999.0, -999.0, 334.38266, 334.4101, 334.43558, 334.45862, 334.4788, 334.49542, 334.50766, 334.51453, 334.51508, 334.50854, 334.49442, 334.47232, 334.44183, 334.40488, 334.35962, 334.30594, 334.24393, 334.17365, 334.09525, 334.00882, 333.91714, 333.8192, 333.71402, 333.6018, 333.48276, 333.36108, 333.23434, -999.0, 332.96356, 332.8252, 332.68317, 332.53748, -999.0, -999.0, 332.10025, 331.95383, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 331.00223, 330.88385, 330.771, 330.66473, 330.56708, 330.47937, 330.39975, 330.32855, 330.26553, 330.21033, 330.1626, 330.1223, 330.0891, 330.06128, 330.0381, 330.0188, 330.00247, 329.98813, 329.97482, 329.96164, 329.9478, 329.93256, -999.0, -999.0, -999.0, 329.84573, 329.81662, 329.78452, 329.74982, 329.7132, 329.6762, 329.63794, 329.5989, 329.55957, 329.52042, 329.48193, 329.44476, 329.40945, 329.37665, 329.34692, 329.322, 329.30096, 329.28424, 329.27222, 329.26474, 329.26358, 329.268, 329.2781, 329.29355, 329.31384, -999.0, 329.36716, 329.3987, 329.4323, 329.4671, 329.50308, -999.0, -999.0, 329.60617, 329.63626, 329.66354, 329.6878, 329.70892, 329.72662, 329.74057, 329.7504, 329.75577, 329.75647, 329.7527, 329.7447, 329.73267, 329.71695, -999.0, -999.0, 329.6508, 329.62363, 329.5953, 329.56732, 329.53894, 329.51074, 329.48325, 329.45706, 329.4327, 329.41107, 329.395, 329.3884, 329.37854, 329.37375, 329.37427, -999.0, -999.0, -999.0, 329.43146, 329.45807, 329.48828, 329.5217, 329.55792, 329.59653, 329.63742, -999.0, -999.0, 329.77237, 329.8181, 329.86328, 329.9074, 329.9501, 329.991, 330.0297, 330.06598, 330.09976, 330.13092, 330.1593, 330.1848, 330.20728, 330.22696, 330.2433, -999.0, 330.2652, 330.27054, 330.2719, 330.26923, 330.26233, 330.2511, -999.0, 330.2156, 330.1922, 330.16586, 330.13712, 330.1067, 330.07526, 330.0436, 330.01297, 329.98428, 329.95654, 329.92984, 329.90427, 329.8797, 329.856, 329.83286, 329.8101, 329.78906, 329.76816, 329.74667, 329.72424, 329.70068, 329.6758, 329.6497, 329.62433, -999.0, -999.0, -999.0, 329.50928, 329.4791, 329.44986, 329.4206, 329.39175, 329.36377, 329.3346, 329.31198, 329.29184, 329.27432, 329.25977, 329.24838, 329.2405, 329.23615, 329.23526, 329.23776, 329.24356, 329.25247, 329.26447, 329.27893, 329.2956, 329.3142, 329.3345, 329.35623, 329.37915, 329.40323, 329.42807, 329.4407, 329.4663, 329.49213, 329.5181, 329.5441, 329.57, 329.59573, 329.62112, 329.646, 329.67023, 329.69363, 329.71603, 329.73724, 329.75702, 329.77524, 329.79184, 329.8068, 329.8201, 329.8317, 329.84174, 329.85022, 329.85727, 329.86295, 329.8674, 329.87076, 329.87314, 329.87466, 329.87558, 329.8761, 329.87646, 329.8769, 329.87772, 329.8795, 329.88208, 329.88583, 329.89105, 329.89813, 329.9074, 329.91922, 329.9336, 329.9505, 329.9699, 329.99176, 330.01584, 330.04202, 330.0695, -999.0, -999.0, -999.0, 330.18912, 330.2217, 330.25558, 330.29095, 330.32794, 330.36667, 330.40698, 330.44876, 330.49176, 330.53586, 330.58194, 330.62848, 330.67517, 330.72168, 330.7678, 330.8133, 330.858, 330.90182, 330.94513, 330.9884, 331.03207, 331.07663, 331.1227, 331.17123, 331.2218, 331.27463, 331.32944, 331.38583, 331.44345, 331.50183, 331.56015, 331.61758, 331.67328, 331.70554, 331.75702, 331.80536, 331.85046, 331.89215, 331.9299, 331.964, 331.99466, 332.0222, 332.0469, 332.06924, 332.08963, 332.1085, -999.0, -999.0, -999.0, 332.17392, 332.18893, 332.20392, 332.2192, 332.23508, 332.25174, 332.2694, 332.28827, 332.30853, 332.3303, 332.35358, 332.37848, 332.40503, 332.43307, 332.46237, 332.4926, 332.52353, 332.55487, 332.58633, 332.61755, 332.64832, 332.6784, 332.70776, 332.73624, 332.76382, 332.79053, 332.8165, 332.84192, 332.86694, 332.89178, 332.91672, 332.94202, 332.96802, 332.9948, 333.02246, 333.051, 333.08044, 333.11072, 333.14154, 333.17273, 333.204, 333.23495, 333.26514, 333.29395, 333.33, 333.35483, 333.37735, 333.3974, 333.41486, 333.4301, 333.4437, 333.45563, 333.46637, 333.4764, 333.48627, 333.4965, 333.5077, 333.52017, 333.53418, 333.54996, 333.5677, 333.5875, 333.60947, 333.6337, 333.66022, 333.68906, 333.7044, 333.73688, 333.77182, 333.8092, 333.84888, 333.8906, 333.93405, 333.97903, 334.0251, 334.07175, 334.12323, 334.16965, 334.21524, 334.25955, 334.3022, 334.34262, 334.38058, 334.41595, 334.44852, 334.47803, 334.50446, 334.5277, 334.54773, 334.56442, 334.57776, 334.5877, 334.59418, 334.59714, 334.5964, 334.59183, 334.58322, 334.57043, 334.55307, 334.5308, 334.5032, 334.4699, 334.4323, 334.3884, 334.33755, 334.2793, 334.21323, 334.13895, 334.0578, 333.96957, 333.87323, 333.76935, -999.0, 333.546, 333.4283, 333.30756, 333.1867, 333.06845, 332.95163, 332.83762, 332.73016, 332.62964, 332.53568, 332.44937, 332.37262, 332.3072, 332.25128, 332.2269, 332.18536, 332.15344, 332.1308, 332.1168, 332.11142, 332.11337, 332.1217, 332.13568, 332.15472, 332.17813, 332.20557, 332.23694, 332.27213, 332.3111, 332.35388, 332.40067, 332.4517, 332.50717, 332.56732, 332.63248, 332.7031, 332.78018, 332.86316, 332.95193, 333.04642, 333.1466, 333.25195, 333.36163, 333.47476, 333.5904, 333.70767, 333.82635, 333.9453, 334.06287, 334.17807, 334.29022, 334.39853, 334.50223, 334.60065, 334.69336, 334.77985, 334.82062, 334.89697, 334.96652, 335.02933, 335.08557, 335.13538, 335.17917, 335.21738, 335.25043, 335.2788, 335.30508, 335.32492, 335.34146, 335.35617, 335.36807, 335.37732, 335.3841, 335.38855, 335.39075, 335.39072, 335.38855, 335.38425, 335.37833, 335.3713, 335.3621, 335.3506, 335.33685, 335.3208, 335.3025, 335.28186, 335.25897, 335.2356, 335.21027, 335.18286, 335.15347, 335.12216, 335.08896, 335.05392, 335.01828, 334.98203, 334.9444, 334.90558, 334.86566, 334.8248, 334.78314, 334.74216, 334.70142, 334.66046, 334.61954, 334.57898, 334.5392, 334.5008, 334.46597, 334.43356, 334.4038, 334.37695, 334.35333, 334.33313, 334.3164, 334.30338, 334.29474, 334.28925, 334.2866, 334.28644, 334.28842, 334.29218, 334.2973, 334.3034, 334.31006, 334.31693, 334.32376, 334.33127, 334.3385, 334.34525, 334.3514, 334.35703, 334.36203, 334.3665, 334.3703, 334.3734, 334.37576, 334.3773, 334.378, 334.379, 334.37927, 334.37885, 334.37787, 334.37643, 334.37476, 334.3729, 334.37097, 334.36902, 334.36716, 334.3654, 334.36417, 334.3637, 334.3635, 334.36353, 334.36386, 334.3646, 334.36575, 334.36737, 334.36835, 334.37057, 334.37317, 334.37607, 334.37918, 334.3824, 334.38577, 334.3896, 334.39316, 334.39648, 334.3998, 334.40247, 334.40472, 334.40662, 334.40808, 334.40912, 334.4097, 334.40985, 334.4096, 334.409, 334.40808, 334.40695, 334.40625, 334.40567, 334.40506, 334.40433, 334.40338, 334.40213, 334.40054, 334.39847, 334.39594, 334.3928, 334.389, 334.38455, 334.37933, 334.37335, 334.36688, 334.36, 334.35208, 334.34308, 334.3329, 334.3215, 334.3088, 334.2948, 334.27942, 334.26266, 334.2446, 334.2252, 334.2053, 334.1844, 334.16226, 334.13898, 334.1146, 334.08926, 334.06305, 334.03613, 334.0086, 333.98062, 333.953, 333.9256, 333.89816, 333.87094, 333.8442, 333.81818, 333.79312, 333.76953, 333.74774, 333.72824, 333.71194, 333.70093, 333.69623, 333.6992, 333.7101, 333.72784, 333.75116, 333.7788, 333.80957, 333.84225, 333.8756, 333.90848, 333.94003, 333.96994, 333.9842, 334.01108, 334.03568, 334.05795, 334.0779, 334.09564, 334.11124, 334.12485, 334.13696, 334.14807, 334.15787, 334.16666, 334.17468, 334.18216, 334.18936, 334.19638, 334.20337, 334.2104, 334.21753, 334.2254, 334.23383, 334.2423, 334.2508, 334.2592, 334.26743, 334.27536, 334.28293, 334.2899, 334.29672, 334.30286, 334.30768, 334.31116, 334.3134, 334.31433, 334.31412, 334.3129, 334.31088, 334.30853, 334.30646, 334.30408, 334.30145, 334.29846, 334.2957, 334.2929, 334.29028, 334.28787, 334.2857, 334.2839, 334.28244, 334.2817, 334.28174, 334.28217, 334.28293, 334.284, 334.28537, 334.28696, 334.28876, 334.29068, 334.2927, 334.2948, 334.29694, 334.2991, 334.30124, 334.3035, 334.30624, 334.30905, 334.31186, 334.31464, 334.3174, 334.3201, 334.32272, 334.32532, 334.32797, 334.3307, 334.33362, 334.33673, 334.34006, 334.3438, 334.3482, 334.3528, 334.3576, 334.36252, 334.36755, 334.37265, 334.3778, 334.383, 334.38818, 334.3933, 334.39838, 334.40332, 334.40866, 334.41403, 334.4192, 334.42404, 334.42862, 334.43283, 334.43668, 334.44016, 334.4432, 334.4458, 334.44824, 334.4508, 334.45288, 334.45453, 334.45587, 334.45697, 334.45795, 334.4589, 334.46005, 334.46152, 334.4644, 334.468, 334.47247, 334.47803, 334.4849, 334.49326, 334.5034, 334.5156, 334.5301, 334.54752, 334.56805, 334.59158, 334.6183, 334.6482, 334.6812, 334.7172, 334.75604, 334.79736, 334.8407, 334.88556, 334.93146, 334.97784, 335.02423, 335.07007, 335.11484, 335.1579, 335.19867, 335.23654, 335.2709, 335.30142, 335.3278, 335.3499, 335.36774, 335.38208, 335.3905, 335.39468, 335.3948, 335.39117, 335.38416, 335.37402, 335.36118, 335.34598, 335.32892, 335.31097, 335.29175, 335.27173, 335.25122, 335.23065, 335.21042, 335.19077, 335.172, 335.15448, 335.13895, 335.1249, 335.1124, 335.10153, 335.09235, 335.08472, 335.0784, 335.07318, 335.06882, 335.06503, 335.0615, 335.0579, 335.05386, 335.04965, 335.04498, 335.0397, 335.03375, 335.02713, 335.01974, 335.01166, 335.0028, 334.9932, 334.98282, 334.9717, 334.95984, 334.94733, 334.9343, 334.9212, 334.9081, 334.89474, 334.88107, 334.8671, 334.8528, 334.83832, 334.82373, 334.80917, 334.79474, 334.78094, 334.76797, 334.75565, 334.7441, 334.73343, 334.72366, 334.71484, 334.70706, 334.70026, 334.69437, 334.68936, 334.68512, 334.6819, 334.67935, 334.67722, 334.67535, 334.67358, 334.67273, 334.67096, 334.669, 334.66678, 334.6642, 334.66135, 334.65808, 334.6544, 334.65036, 334.64627, 334.6442, 334.6398, 334.63516, 334.6305, 334.6259, 334.62152, 334.6175, 334.61392, 334.61087, 334.60843, 334.60648, 334.60532, 334.60516, 334.60553, 334.6064, 334.60782, 334.60974, 334.6122, 334.6153, 334.619, 334.6234, 334.62857, 334.6345, 334.64117, 334.64865, 334.65695, 334.66592, 334.6755, 334.68555, 334.69595, 334.7012, 334.71164, 334.7217, 334.7311, 334.7395, 334.7464, 334.7513, 334.75406, 334.75397, 334.75058, 334.74347, 334.73837, 334.72488, 334.7069, 334.68445, 334.6575, 334.62604, 334.5904, 334.5509, 334.50793, 334.4622, 334.41434, 334.3897, 334.33945, 334.28848, 334.23746, 334.1871, 334.1381, 334.0912, 334.047, 334.00616, 333.96933, 333.93716, 333.9104, 333.88934, 333.87454, 333.86655, 333.86618, 333.87476, 333.89362, 333.92407, 333.96634, 334.01877, 334.0795, 334.14667, 334.21838, 334.29227, 334.36575, 334.43652, 334.50272, 334.56375, 334.61908, 334.66815, 334.71066, 334.7468, 334.77676, 334.80078, 334.81918, 334.83255, 334.84143, 334.84653, 334.84842, 334.84763, 334.84467, 334.84256, 334.83746, 334.83157, 334.8253, 334.81912, 334.8135, 334.8087, 334.80487, 334.80228, 334.80112, 334.80112, 334.8024, 334.80554, 334.81064, 334.81778, 334.82697, 334.83807, 334.8511, -999.0, -999.0, -999.0, -999.0, 334.93185, 334.95428, 334.9781, 335.0031, 335.02924, 335.05634, 335.08438, 335.11322, 335.1279, 335.15784, 335.17615, 335.20715, 335.2389, 335.27124, 335.3041, 335.3373, 335.3707, 335.40405, 335.43713, 335.4699, 335.5018, 335.5325, 335.562, 335.59036, 335.6176, 335.64386, 335.66922, 335.69373, 335.71753, 335.7407, 335.7634, 335.78586, 335.8082, 335.83063, 335.85333, 335.87653, 335.90045, 335.92523, 335.95114, 335.9783, 336.00696, 336.0219, 336.05307, 336.08597, 336.12064, 336.1571, 336.19534, 336.2353, 336.27682, 336.31982, 336.36417, 336.4097, 336.45578, 336.502, 336.54788, 336.59277, 336.636, 336.67682, 336.71463, 336.74893, 336.77914, 336.80478, 336.82553, 336.84146, 336.8527, 336.85938, 336.86185, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 338.65753, 338.68747, 338.7102, 338.72485, 338.7305, 338.72626, 338.71207, 338.68964, 338.66092, 338.62778, 338.59183, 338.5541, 338.51556, 338.4772, 338.43982, 338.40402, 338.37048, 338.33923, 338.3106, 338.2846, 338.26126, 338.24057, 338.22247, 338.2069, 338.19366, 338.18265, 338.17368, 338.1665, 338.16104, 338.15732, 338.15472, 338.15295, 338.15167, 338.1506, 338.1494, 338.1479, 338.14575, 338.14282, 338.1388, 338.13354, 338.1268, 338.11853, 338.11392, 338.10333, 338.0911, 338.07724, 338.06192, 338.04526, 338.0275, 338.0088, 337.9894, 337.96942, 337.94916, 337.92905, 337.9087, 337.8882, 337.86765, 337.84708, 337.82657, 337.8061, 337.78555, 337.7649, 337.74405, 337.7337, 337.71326, 337.69287, 337.67267, 337.6528, 337.6335, 337.61502, 337.59756, 337.58133, 337.56647, 337.55304, 337.54117, 337.5311, 337.52283, 337.51608, 337.51074, 337.50674, 337.50394, 337.50208, 337.501, 337.50055, 337.5006, 337.5012, 337.50217, 337.50354, 337.5053, 337.50754, 337.51022, 337.51352, 337.5176, 337.52274, 337.52805, 337.53394, 337.54037, 337.5472, 337.55438, 337.56177, 337.56924, 337.57675, 337.58414, 337.59137, 337.59845, 337.6054, 337.61224, 337.61902, 337.6257, 337.63226, 337.6387, 337.645, 337.65118, 337.65747, 337.66373, 337.6668, 337.67294, 337.67896, 337.6848, 337.69055, 337.69608, 337.70135, 337.70633, 337.7109, 337.7151, 337.71878, 337.72195, 337.72458, 337.72662, 337.72815, 337.72916, 337.72968, 337.72974, 337.72943, 337.72876, 337.7278, 337.72684, 337.7258, 337.72464, -999.0, -999.0, 337.7214, 337.72104, 337.7213, 337.7224, 337.7244, 337.7273, 337.72913, 337.73355, 337.73886, -999.0, -999.0, -999.0, -999.0, -999.0, 337.7838, 337.78775, 337.7951, 337.80154, 337.8067, 337.81024, 337.81195, 337.81174, 337.80945, 337.80508, 337.79855, 337.78998, 337.7849, 337.77368, 337.76062, 337.7456, 337.72864, 337.70972, 337.68884, 337.66647, 337.643, 337.6189, 337.59464, 337.58264, 337.55945, 337.5381, 337.5189, 337.50266, 337.49033, 337.4828, 337.48096, 337.48523, -999.0, 337.51462, 337.5384, 337.5673, 337.5995, 337.63306, 337.6664, 337.6985, 337.7288, 337.75677, 337.78204, 337.80444, 337.81458, 337.83267, 337.84793, 337.86044, 337.8705, 337.87854, 337.88486, 337.88977, 337.8938, 337.8969, 337.89914, 337.9, 337.90112, 337.9014, 337.9008, 337.89917, 337.89655, 337.89285, 337.88806, 337.88266, 337.87613, 337.86853, 337.86432, 337.8551, 337.84485, 337.83356, 337.8212, 337.80783, 337.7936, 337.77866, 337.7627, 337.74567, 337.73676, 337.7181, 337.69824, 337.67703, 337.65442, 337.63095, 337.60645, 337.58102, 337.55493, 337.5285, 337.5022, 337.4764, 337.45212, 337.4298, 337.41055, 337.3955, 337.3858, 337.38187, 337.38373, 337.39142, 337.40506, 337.4138, 337.43427, 337.4577, 337.48282, 337.50854, 337.53458, 337.5606, 337.58646, 337.61188, 337.63684, 337.66162, 337.68585, 337.7095, 337.7328, 337.7558, 337.7787, 337.80164, 337.82465, 337.84772, 337.87094, 337.89423, 337.9175, 337.94064, 337.96353, 337.9861, 338.0081, 338.02924, 338.04932, 338.06818, 338.08554, 338.10117, 338.10822, 338.1207, 338.1309, 338.13882, 338.1445, 338.14786, 338.14908, 338.14832, 338.14597, 338.14203, 338.13953, 338.13358, 338.12653, 338.11862, 338.11005, 338.101, 338.09167, 338.08218, 338.07272, 338.06342, 338.05365, 338.0455, 338.038, 338.0313, 338.02563, 338.02118, 338.01807, 338.01642, 338.01633, 338.01785, 338.0211, 338.02332, 338.02908, 338.0365, 338.04556, 338.05618, 338.06833, 338.08188, 338.09677, 338.11288, 338.13013, 338.14856, 338.1581, 338.17795, 338.1988, 338.22076, 338.24396, 338.26846, 338.2945, 338.32224, 338.3519, 338.3836, 338.41745, 338.43518, 338.47226, 338.51157, 338.5529, 338.59595, 338.64047, 338.68613, 338.73248, 338.77908, 338.82538, 338.87085, 338.8932, 338.93683, 338.9789, 339.01923, 339.05753, 339.09384, 339.1282, 339.1607, 339.19135, 339.22018, 339.24738, 339.26035, 339.28497, 339.30783, 339.32883, 339.34784, 339.36484, 339.37964, 339.39212, 339.40216, 339.4096, 339.4144, 339.41653, 339.416, 339.41287, 339.4074, 339.3996, 339.38968, 339.37787, 339.3644, 339.34967, 339.33398, 339.31772, 339.3012, 339.28503, 339.2698, 339.25592, 339.24377, 339.23376, 339.22644, 339.22217, 339.22122, 339.22202, 339.22604, 339.23337, 339.24396, 339.25748, 339.2736, 339.29193, 339.3121, 339.33386, 339.35907, 339.3827, 339.4066, 339.4305, 339.45416, 339.47726, 339.49957, 339.5211, 339.54175, 339.56155, 339.58047, 339.58963, 339.60724, 339.62405, 339.64005, 339.65524, 339.66968, 339.68338, 339.69635, 339.70856, 339.7201, 339.7309, 339.74088, 339.74997, 339.75812, 339.76517, 339.77112, 339.77594, 339.77975, 339.7827, 339.78488, 339.78644, 339.78705, 339.788, 339.78873, 339.78946, 339.7903, 339.7915, 339.7933, 339.7957, 339.79874, 339.80258, 339.80478, 339.80988, 339.8159, 339.82278, 339.83066, 339.83948, 339.8493, 339.8601, 339.87198, 339.88492, 339.89883, 339.91367, 339.92133, -999.0, 339.95355, 339.97034, 339.9874, 340.00446, 340.02142, 340.03818, 340.0547, 340.07083, 340.08655, 340.10184, 340.11664, 340.1309, 340.14462, 340.1579, 340.17078, 340.18338, 340.19583, 340.2082, 340.2144, 340.22687, 340.2396, 340.25256, 340.26596, 340.2796, 340.2935, 340.30753, 340.32147, 340.33517, -999.0, 340.36118, 340.36737, 340.3794, 340.391, 340.40225, 340.41318, 340.42386, 340.4343, 340.44458, 340.45468, 340.4645, 340.47418, 340.48352, 340.49243, -999.0, -999.0, -999.0, -999.0, 340.52887, 340.53433, 340.53918, 340.5418, 340.5458, 340.5493, 340.55237, 340.555, 340.55704, 340.5584, 340.55914, 340.55893, 340.5576, 340.55646, 340.55316, 340.54834, 340.54196, 340.534, 340.52438, 340.51315, 340.5004, 340.48627, 340.4709, 340.45447, 340.43713, 340.41895, 340.39996, 340.38034, -999.0, -999.0, -999.0, -999.0, -999.0, 340.2685, 340.25876, 340.23987, 340.2217, -999.0, -999.0, -999.0, 340.15887, 340.14642, -999.0, -999.0, 340.1191, 340.11407, 340.11154, 340.11182, 340.11554, 340.12344, 340.1363, 340.15488, -999.0, 340.20828, 340.2414, 340.2776, 340.31613, 340.35632, 340.39743, 340.4388, 340.48004, 340.52097, 340.56146, 340.60135, 340.64062, 340.6794, 340.7178, 340.73688, 340.77487, 340.81268, 340.85037, 340.88806}
theta_v =
  {313.1811, -999.0, -999.0, -999.0, -999.0, -999.0, 313.2171, 313.21448, 313.2115, 313.20798, 313.20398, 313.19952, 313.1946, 313.18927, 313.18356, 313.17755, 313.1714, 313.1651, 313.15894, 313.15314, 313.14795, 313.14355, 313.1402, 313.13803, 313.1373, 313.13812, 313.14062, 313.1449, 313.15097, 313.1589, 313.16858, 313.17975, 313.19226, 313.2059, 313.2204, 313.23553, 313.25107, 313.2667, 313.2823, 313.29767, 313.31268, 313.32715, 313.34094, 313.354, 313.36624, 313.3776, 313.38812, 313.39798, 313.40723, 313.41605, 313.42453, 313.43283, 313.44107, 313.44946, 313.45825, 313.4677, -999.0, 313.4899, 313.50336, 313.51892, 313.53897, 313.56027, 313.58475, 313.61258, 313.644, 313.67914, 313.71808, 313.76083, 313.80743, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 314.52026, -999.0, -999.0, -999.0, 314.71225, 314.7528, 314.7897, 314.8222, 314.84952, 314.871, 314.88666, 314.8965, -999.0, -999.0, -999.0, -999.0, -999.0, 314.85577, 314.83932, 314.82193, 314.80405, 314.78622, 314.7689, 314.7524, -999.0, 314.72345, 314.71143, 314.70096, 314.69214, 314.68484, 314.6789, 314.67407, 314.67007, 314.6667, -999.0, -999.0, 314.65952, 314.6579, 314.6564, 314.65488, 314.6531, 314.6509, 314.6483, 314.64532, 314.64203, 314.63852, 314.63495, 314.63153, 314.62848, 314.62598, 314.62415, 314.62305, 314.62274, 314.6233, 314.6247, 314.6269, 314.6299, 314.63364, 314.638, 314.64276, 314.6478, 314.6529, 314.6579, 314.66266, 314.667, 314.67084, 314.67407, 314.67676, 314.67883, 314.68036, 314.68137, 314.682, 314.68237, 314.68256, 314.68265, 314.68268, 314.68277, 314.68292, 314.68317, 314.68353, 314.68396, 314.68445, 314.68497, 314.68552, 314.6861, 314.6867, 314.68732, 314.68802, 314.6888, 314.68976, 314.6908, 314.69193, 314.69308, 314.69427, 314.69543, 314.69662, 314.69778, 314.69894, 314.7001, 314.70123, 314.70236, 314.70343, 314.70438, 314.70514, 314.7056, 314.7057, 314.70532, 314.70444, 314.70294, 314.70078, 314.69797, 314.69458, 314.6907, 314.68634, 314.68158, 314.6765, 314.67126, 314.66586, 314.66055, 314.65558, 314.65118, 314.64755, 314.64474, 314.6427, 314.64142, 314.6409, 314.64114, 314.64224, 314.64423, 314.64716, 314.65094, 314.65536, 314.66034, 314.6657, 314.6713, 314.677, 314.68262, 314.68808, 314.6934, 314.69864, 314.70386, 314.70914, 314.7147, 314.72073, 314.72754, 314.7353, 314.74405, 314.75385, 314.76474, 314.77673, 314.78964, 314.8033, 314.81754, 314.83212, 314.84683, 314.86142, 314.87564, 314.8893, 314.9022, 314.91415, 314.92502, 314.9346, 314.9429, 314.94986, 314.9555, 314.9598, 314.96283, 314.96457, 314.96506, 314.9644, 314.96262, 314.9599, 314.9564, 314.95218, 314.94742, 314.9423, 314.93695, 314.93155, 314.92627, 314.9212, 314.9165, 314.91235, 314.90887, 314.906, 314.90442, 314.90396, 314.90472, 314.90668, 314.9099, 314.9144, 314.92004, 314.9267, 314.9342, 314.94244, 314.9512, 314.96033, 314.96964, 314.97894, 314.9882, 314.99728, 315.0062, -999.0, -999.0, 315.0312, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 314.7247, 314.71417, 314.70294, 314.69086, 314.67648, 314.66238, 314.64728, 314.63113, 314.61395, 314.596, 314.5776, 314.55905, 314.54065, 314.52267, 314.5054, 314.48904, -999.0, -999.0, 314.44708, 314.43546, 314.42505, 314.41592, -999.0, -999.0, -999.0, -999.0, 314.39398, 314.394, 314.3951, 314.39688, 314.39893, 314.40082, 314.40213, 314.40256, 314.40176, 314.39938, 314.39517, 314.38907, 314.3811, 314.3713, 314.35977, 314.34677, 314.3328, 314.31824, 314.30356, 314.2893, 314.2761, 314.26453, 314.2552, 314.24835, 314.2443, 314.24313, 314.24515, 314.2503, 314.25867, 314.2702, 314.28485, 314.30237, 314.32233, 314.3443, 314.3679, 314.39267, 314.41806, 314.4436, 314.46884, 314.49338, 314.517, 314.53943, 314.56042, 314.57974, 314.59726, 314.61273, 314.62604, 314.637, 314.64554, 314.65155, 314.6549, 314.65558, 314.6535, 314.64862, 314.64093, 314.63043, 314.61722, 314.60135, 314.58292, 314.56207, 314.53903, 314.51404, 314.48724, 314.45898, 314.42953, 314.39923, 314.36838, 314.3376, 314.30743, 314.27863, -999.0, -999.0, 314.20355, 314.18542, 314.1709, 314.15994, 314.1523, 314.1479, 314.14645, 314.1476, 314.15103, 314.1563, 314.16302, 314.171, 314.17993, 314.1896, 314.19983, 314.21045, 314.22137, 314.23245, 314.2436, 314.25476, 314.2659, 314.27707, 314.28815, 314.2992, 314.31018, 314.3211, 314.33194, 314.34268, 314.35324, 314.36356, 314.37357, 314.38324, -999.0, -999.0, 314.409, 314.41623, 314.42267, 314.42825, 314.43286, 314.43655, 314.43927, 314.44104, 314.44183, 314.44168, 314.4407, 314.4389, 314.43637, 314.43317, 314.42938, 314.4251, 314.42047, 314.4155, 314.4103, 314.40497, 314.39954, 314.39407, 314.38858, 314.38306, 314.3775, 314.37195, 314.3664, 314.3608, 314.3553, 314.34985, 314.3446, 314.33966, 314.33514, 314.33118, 314.32788, 314.3255, 314.32413, 314.32388, 314.3249, 314.32727, 314.3311, 314.3365, 314.3437, 314.35278, 314.36395, 314.37735, 314.39316, 314.41153, 314.43262, 314.4565, 314.4833, 314.51303, -999.0, -999.0, 314.62024, 314.66193, -999.0, -999.0, -999.0, -999.0, -999.0, 314.96854, 315.02682, -999.0, -999.0, 315.20468, 315.26318, 315.32043, -999.0, -999.0, 315.48062, -999.0, 315.5753, 315.6186, 315.65927, 315.69748, 315.7367, 315.77, 315.80118, 315.8304, 315.85782, 315.8834, 315.90707, 315.9288, 315.94852, 315.966, 315.9811, 315.9936, -999.0, -999.0, -999.0, 316.0161, 316.0153, 316.01224, 316.00717, 316.00034, 315.99197, 315.98236, 315.97168, 315.9602, 315.9482, 315.9359, 315.92365, 315.91165, 315.9002, 315.88953, 315.87973, 315.87097, 315.86337, 315.857, 315.85184, 315.8479, 315.84518, 315.8436, 315.84302, 315.84332, 315.84436, 315.84604, 315.84824, 315.85086, 315.85382, 315.857, -999.0, -999.0, -999.0, 315.87186, 315.87595, 315.88022, 315.88464, 315.8892, 315.8939, 315.89874, 315.90372, 315.9088, 315.91388, 315.91882, 315.92355, 315.92798, 315.932, 315.93558, -999.0, -999.0, 315.94302, 315.94434, 315.9451, 315.94525, 315.9449, 315.94397, 315.9426, 315.94064, 315.93802, 315.93466, 315.93045, 315.9253, 315.9191, -999.0, 315.90317, 315.89334, 315.88235, 315.87024, 315.85706, 315.8429, 315.82794, 315.81238, 315.79633, 315.77988, 315.76306, 315.74597, 315.72687, 315.7093, 315.6916, 315.67383, 315.65607, 315.63834, 315.6207, 315.6032, 315.5859, 315.56894, 315.55243, 315.53653, 315.5214, 315.5071, 315.49377, 315.48148, 315.47025, 315.46002, 315.45056, 315.44168, 315.4332, 315.42474, 315.41605, 315.4067, 315.39648, 315.38544, 315.37378, 315.36185, 315.34985, 315.3381, 315.32684, 315.3164, 315.307, 315.29877, 315.29156, 315.28537, 315.2801, 315.27545, 315.27097, 315.26624, 315.26083, 315.25452, 315.24716, 315.2387, 315.229, 315.21802, 315.20578, 315.19223, 315.1774, 315.16153, 315.145, 315.12808, 315.1112, 315.09467, 315.07877, 315.06387, 315.05032, 315.0384, 315.02838, 315.02057, 315.01526, 315.01273, 315.0133, 315.0173, 315.02496, 315.03644, 315.05185, 315.07123, 315.0946, 315.1214, 315.1508, 315.18185, 315.21378, 315.24588, 315.27762, 315.3085, 315.338, 315.36618, 315.39337, 315.41992, 315.4462, 315.4726, 315.4995, 315.5274, 315.55658, 315.5871, 315.61874, 315.65137, 315.68472, 315.7184, 315.75198, 315.78497, 315.8169, 315.84763, 315.8772, 315.90567, 315.93307, 315.95947, 315.98492, 316.00946, 316.03314, 316.05606, 316.08054, 316.10217, 316.12332, 316.14398, 316.16412, 316.1837, 316.20264, 316.22086, 316.23837, 316.2551, 316.27103, 316.28607, 316.3003, 316.3137, 316.32623, 316.33795, 316.34882, 316.3588, 316.36792, 316.3762, 316.38373, 316.39056, 316.3968, 316.40256, 316.40802, 316.4133, 316.4186, 316.424, 316.4297, 316.43576, 316.44235, 316.44952, 316.45737, 316.46594, 316.47528, 316.48538, 316.49622, 316.5078, 316.52005, 316.5329, 316.54626, 316.56003, 316.57407, 316.58826, 316.60248, 316.61652, 316.63025, 316.64352, 316.65628, 316.6683, 316.67953, 316.68997, 316.69492, 316.70425, 316.71298, 316.72113, 316.72882, 316.73618, 316.74332, 316.7503, 316.7573, 316.7643, 316.77142, 316.77875, 316.7863, 316.79407, 316.8022, 316.81055, 316.81915, 316.82788, 316.8366, 316.84525, 316.8537, 316.86188, 316.86966, 316.87692, 316.88358, 316.88956, 316.89474, 316.8991, 316.9027, 316.90564, 316.908, 316.90985, 316.91135, 316.91257, -999.0, -999.0, 316.91577, 316.9172, 316.91916, 316.92178, 316.9253, 316.92987, 316.93573, 316.94305, 316.95197, 316.96252, 316.97488, 316.98904, 317.00504, 317.02274, 317.0441, 317.0652, 317.08777, 317.11182, 317.13718, 317.16385, 317.19177, 317.22086, 317.25107, 317.28238, 317.31482, 317.3484, 317.38312, 317.419, -999.0, -999.0, 317.532, 317.57086, 317.60977, 317.64832, 317.686, 317.72247, 317.7573, 317.79007, 317.82043, 317.84808, 317.8729, 317.8948, 317.91376, 317.92975, 317.94296, 317.95358, 317.96188, 317.96808, 317.9725, 317.97543, 317.97723, 317.97818, 317.97858, 317.9787, 317.97885, 317.97922, 317.97998, -999.0, 317.98297, 317.98535, 317.9884, 317.99203, -999.0, -999.0, 318.00595, 318.0109, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 318.0219, 318.01834, 318.01364, 318.00806, 318.00177, 317.99506, 317.98813, 317.98123, 317.97446, 317.9679, 317.9616, 317.9557, 317.95013, 317.94504, 317.94043, 317.9363, 317.93265, 317.9294, 317.9265, 317.92392, 317.92157, 317.91943, -999.0, -999.0, -999.0, 317.91193, 317.9103, 317.90884, 317.9075, 317.90637, 317.90546, 317.9048, 317.90433, 317.90408, 317.904, 317.90405, 317.9043, 317.90475, 317.90543, 317.9064, 317.90768, 317.9093, 317.91135, 317.91382, 317.91693, 317.92007, 317.92346, 317.92697, 317.93054, 317.93405, -999.0, 317.94046, 317.94324, 317.94562, 317.94754, 317.94897, -999.0, -999.0, 317.94965, 317.94852, 317.9467, 317.94427, 317.9413, 317.93787, 317.93414, 317.93027, 317.92645, 317.9229, 317.91992, 317.9179, 317.91714, 317.91797, -999.0, -999.0, 317.93265, 317.94247, 317.95514, 317.97086, 317.98978, 318.01212, 318.03802, 318.06763, 318.101, 318.1383, 318.17953, 318.20166, 318.24884, 318.30002, 318.355, -999.0, -999.0, -999.0, 318.60806, 318.67804, 318.74997, 318.82343, 318.89804, 318.97333, 319.04895, -999.0, -999.0, 319.2727, 319.34442, 319.41373, 319.4801, 319.54306, 319.6021, 319.6568, 319.70688, 319.75232, 319.7931, 319.8292, 319.86075, 319.888, 319.91122, 319.9307, -999.0, 319.95953, 319.9695, 319.977, 319.98227, 319.98566, 319.98746, -999.0, 319.98767, 319.98682, 319.98587, 319.98526, 319.9853, 319.98633, 319.98865, 319.99258, 319.99832, 320.00592, 320.01553, 320.0272, 320.04095, 320.05667, 320.07428, 320.09372, 320.1148, 320.13733, 320.16113, 320.186, 320.2118, 320.23834, 320.26556, 320.2933, -999.0, -999.0, -999.0, 320.40656, 320.43457, 320.4621, 320.48886, 320.5147, 320.5395, 320.56546, 320.58783, 320.60895, 320.62888, 320.64767, 320.66544, 320.68216, 320.698, 320.71298, 320.7272, 320.74075, 320.75372, 320.7662, 320.7783, 320.79013, 320.8018, 320.81332, 320.8248, 320.83633, 320.8479, 320.85956, 320.8654, 320.87714, 320.88898, 320.90085, 320.91272, 320.92453, 320.93628, 320.94788, 320.95926, 320.9703, 320.981, 320.99127, 321.00113, 321.0105, 321.0194, 321.02783, 321.03586, 321.0435, 321.05075, 321.05768, 321.06436, 321.0708, 321.07706, 321.0832, 321.08923, 321.09525, 321.10123, 321.10724, 321.11325, 321.11932, 321.12543, 321.13153, 321.13757, 321.14355, 321.1494, 321.1552, 321.16092, 321.16663, 321.17233, 321.17807, 321.18387, 321.18976, 321.19577, 321.20184, 321.20798, 321.21408, -999.0, -999.0, -999.0, 321.23868, 321.24503, 321.25156, 321.25836, 321.26544, 321.2729, 321.28076, 321.28903, 321.2978, 321.307, 321.31665, 321.3267, 321.33707, 321.34772, 321.35864, 321.3698, 321.38116, 321.3927, 321.40454, 321.41672, 321.4294, 321.4427, 321.4567, 321.47156, 321.4874, 321.5043, 321.52225, 321.54117, 321.561, 321.5817, 321.60297, 321.62463, 321.64642, 321.65942, 321.68094, 321.70206, 321.72256, 321.74234, 321.76126, 321.77927, 321.79623, 321.81213, 321.8269, 321.84045, 321.85278, 321.8638, -999.0, -999.0, -999.0, 321.8965, 321.90244, 321.90784, 321.91296, 321.91806, 321.9233, 321.92886, 321.93497, 321.9417, 321.94922, 321.95752, 321.96664, 321.97665, 321.98755, 321.9994, 322.01215, 322.02588, 322.0406, 322.05634, 322.07312, 322.09094, 322.1098, 322.12964, 322.15045, 322.17212, 322.19467, 322.21805, 322.24228, 322.2673, 322.29318, 322.31998, 322.3477, 322.37643, 322.40613, 322.43677, 322.46826, 322.5005, 322.5334, 322.56677, 322.6005, 322.63437, 322.66815, 322.70148, 322.73398, 322.7741, 322.80405, 322.8324, 322.859, 322.8837, 322.90652, 322.92764, 322.94724, 322.96548, 322.9826, 322.99872, 323.01404, 323.02875, 323.043, 323.05698, 323.07086, 323.08478, 323.09897, 323.11365, 323.129, 323.1453, 323.16272, 323.1719, 323.1914, 323.21252, 323.2354, 323.2601, 323.2865, 323.31458, 323.34427, 323.37534, 323.4075, 323.44388, 323.47757, 323.5115, 323.5454, 323.57895, 323.61188, 323.64398, 323.67508, 323.70505, 323.73367, 323.76096, 323.78674, 323.81107, 323.8338, 323.85498, 323.87466, 323.89285, 323.90958, 323.92487, 323.93875, 323.9513, 323.96252, 323.97238, 323.9808, 323.98773, 323.99307, 323.99673, 323.9985, 323.99823, 323.9957, 323.99078, 323.98328, 323.973, 323.95984, 323.94388, 323.9253, -999.0, 323.88113, 323.85632, 323.8304, 323.80402, 323.7777, 323.75204, 323.72757, 323.70486, 323.68445, 323.66666, 323.65192, 323.64053, 323.63287, 323.62888, 323.62827, 323.6298, 323.6349, 323.6434, 323.65506, 323.66953, 323.68652, 323.7057, 323.72678, 323.7495, 323.77356, 323.7988, 323.82523, 323.8529, 323.88177, 323.91196, 323.9437, 323.97708, 324.0124, 324.04984, 324.08966, 324.13214, 324.17755, 324.2261, 324.27786, 324.33292, 324.39142, 324.45328, 324.51813, 324.5857, 324.6557, 324.72775, 324.80142, 324.87625, 324.95187, 325.0278, 325.10364, 325.17892, 325.25333, 325.32635, 325.39774, 325.46707, 325.5009, 325.56662, 325.62976, 325.69028, 325.74814, 325.8033, 325.85593, 325.90613, 325.95407, 325.99988, 326.04797, 326.08972, 326.1297, 326.16803, 326.20474, 326.2399, 326.27353, 326.3057, 326.33633, 326.36554, 326.39325, 326.41953, 326.4443, 326.46762, 326.48944, 326.5098, 326.5287, 326.5461, 326.56213, 326.5768, 326.59012, 326.6021, 326.61285, 326.62234, 326.6306, 326.6377, 326.64365, 326.64844, 326.65222, 326.65503, 326.65698, 326.65817, 326.6587, 326.65866, 326.65814, 326.65726, 326.6562, 326.65512, 326.6542, 326.65372, 326.65387, 326.65494, 326.65723, 326.66098, 326.66632, 326.6734, 326.68228, 326.69308, 326.70572, 326.72015, 326.73627, 326.754, 326.7732, 326.7936, 326.8151, 326.83746, 326.86053, 326.8841, 326.90796, 326.93195, 326.956, 326.98, 327.0039, 327.02765, 327.05115, 327.07446, 327.0975, 327.12027, 327.1427, 327.1647, 327.18622, 327.20718, 327.2276, 327.2474, 327.26663, 327.28528, 327.3034, 327.3211, 327.33847, 327.35562, 327.37256, 327.38937, 327.4061, 327.42276, 327.4394, 327.45602, 327.47266, 327.48932, 327.50607, 327.5229, 327.53986, 327.55695, 327.56555, 327.5828, 327.60013, 327.61746, 327.6348, 327.65204, 327.66913, 327.686, 327.7026, 327.7189, 327.73648, 327.75208, 327.7673, 327.78217, 327.79663, 327.81073, 327.82446, 327.8379, 327.85098, 327.86383, 327.87646, 327.88898, 327.9014, 327.91382, 327.92624, 327.9387, 327.95105, 327.96335, 327.97552, 327.98755, 327.99936, 328.01096, 328.02225, 328.03323, 328.04385, 328.05405, 328.06378, 328.07294, 328.0815, 328.0894, 328.09653, 328.10284, 328.10834, 328.11295, 328.11664, 328.11945, 328.12134, 328.12238, 328.1226, 328.12195, 328.1205, 328.1183, 328.1153, 328.1116, 328.10724, 328.1023, 328.0968, 328.09085, 328.08453, 328.0779, 328.07117, 328.0644, 328.0578, 328.05154, 328.04584, 328.04105, 328.03745, 328.0354, 328.0356, 328.0392, 328.0474, 328.06125, 328.08112, 328.10608, 328.13525, 328.1677, 328.2025, 328.23883, 328.27573, 328.31232, 328.348, 328.3826, 328.39944, 328.4321, 328.46326, 328.49298, 328.52136, 328.5485, 328.57455, 328.59964, 328.624, 328.6478, 328.6712, 328.69446, 328.7177, 328.7412, 328.76514, 328.78955, 328.8145, 328.84006, 328.86627, 328.893, 328.92023, 328.9478, 328.97562, 329.00354, 329.03146, 329.05917, 329.08655, 329.11334, 329.1393, 329.16418, 329.18774, 329.2099, 329.23062, 329.24994, 329.26782, 329.28442, 329.2999, 329.31442, 329.3282, 329.34125, 329.35376, 329.36697, 329.3786, 329.38992, 329.40106, 329.4121, 329.42316, 329.43423, 329.4454, 329.45676, 329.46826, 329.47998, 329.4919, 329.50397, 329.51624, 329.52863, 329.54117, 329.55386, 329.56668, 329.5796, 329.59262, 329.60574, 329.61896, 329.63226, 329.64566, 329.65918, 329.6728, 329.6865, 329.70026, 329.71402, 329.72775, 329.74155, 329.75537, 329.76935, 329.7835, 329.79788, 329.81244, 329.8273, 329.84238, 329.8578, 329.87344, 329.88943, 329.90573, 329.92236, 329.9393, 329.95654, 329.97412, 329.992, 330.01016, 330.0285, 330.04706, 330.06573, 330.0845, 330.1033, 330.12207, 330.1408, 330.15942, 330.17792, 330.19623, 330.21436, 330.23227, 330.24994, 330.26736, 330.2846, 330.30173, 330.3188, 330.3359, 330.35318, 330.37076, 330.3888, 330.40744, 330.42682, 330.44705, 330.46832, 330.49072, 330.51437, 330.5394, 330.56595, 330.59415, 330.6241, 330.65594, 330.68973, 330.72556, 330.76337, 330.80304, 330.84448, 330.88754, 330.93195, 330.97736, 331.02353, 331.07007, 331.11667, 331.16302, 331.20874, 331.2535, 331.2969, 331.3385, 331.3779, 331.41464, 331.44852, 331.4793, 331.50684, 331.53094, 331.55356, 331.5707, 331.58475, 331.59583, 331.60413, 331.60995, 331.61353, 331.61508, 331.6149, 331.61325, 331.61035, 331.6065, 331.60196, 331.597, 331.59186, 331.58688, 331.58224, 331.5781, 331.57465, 331.57205, 331.57037, 331.56973, 331.5701, 331.5716, 331.574, 331.57724, 331.58105, 331.58533, 331.5898, 331.59427, 331.59848, 331.6022, 331.60544, 331.60815, 331.6104, 331.61218, 331.61356, 331.61453, 331.6152, 331.61557, 331.6157, 331.61557, 331.61523, 331.61462, 331.61386, 331.61298, 331.61203, 331.6111, 331.61017, 331.6092, 331.6081, 331.60687, 331.60553, 331.6042, 331.6028, 331.60156, 331.60046, 331.5996, 331.59912, 331.5991, 331.59955, 331.60056, 331.60214, 331.60434, 331.60715, 331.61053, 331.61453, 331.6191, 331.62415, 331.62964, 331.63547, 331.64157, 331.64786, 331.65103, 331.65747, 331.66388, 331.67026, 331.6765, 331.6826, 331.68842, 331.69403, 331.69934, 331.7044, 331.70682, 331.71146, 331.71594, 331.72043, 331.72504, 331.7299, 331.73514, 331.7408, 331.74698, 331.7537, 331.7617, 331.7694, 331.7775, 331.78583, 331.79443, 331.8032, 331.81204, 331.821, 331.83008, 331.83923, 331.84854, 331.85803, 331.86774, 331.87772, 331.88803, 331.89874, 331.90982, 331.9213, 331.93314, 331.94534, 331.9515, 331.9639, 331.97617, 331.98813, 331.99948, 332.00992, 332.01898, 332.0264, 332.0317, 332.03455, 332.0345, 332.03323, 332.02814, 332.01944, 332.00702, 331.9908, 331.97076, 331.94705, 331.91992, 331.8896, 331.85638, 331.82074, 331.8022, 331.76398, 331.7247, 331.68497, 331.64536, 331.60654, 331.5691, 331.5336, 331.5007, 331.47095, 331.44492, 331.42325, 331.4064, 331.39496, 331.38943, 331.39062, 331.39975, 331.41797, 331.44656, 331.48572, 331.534, 331.58984, 331.65167, 331.71774, 331.78592, 331.85413, 331.92023, 331.98267, 332.04083, 332.09415, 332.1421, 332.18436, 332.221, 332.25214, 332.27792, 332.29852, 332.31445, 332.32617, 332.3341, 332.33878, 332.34067, 332.34024, 332.33932, 332.3364, 332.33234, 332.32755, 332.32248, 332.31754, 332.31296, 332.30896, 332.30573, 332.30347, 332.30276, 332.30228, 332.30313, 332.30554, 332.30957, 332.3152, 332.3224, 332.33112, -999.0, -999.0, -999.0, -999.0, 332.38858, 332.4051, 332.42273, 332.44147, 332.46118, 332.48178, 332.50317, 332.5253, 332.53662, 332.5597, 332.57385, 332.59787, 332.62253, 332.6477, 332.67337, 332.69934, 332.72552, 332.75177, 332.77786, 332.80356, 332.8286, 332.8528, 332.87616, 332.89868, 332.92044, 332.94153, 332.962, 332.98193, 333.0014, 333.0205, 333.03934, 333.0581, 333.07693, 333.096, 333.11548, 333.1355, 333.15622, 333.17783, 333.20044, 333.22418, 333.24918, 333.26218, 333.28925, 333.31775, 333.34766, 333.37903, 333.41183, 333.44598, 333.4814, 333.5181, 333.55582, 333.59436, 333.63336, 333.67255, 333.71152, 333.74976, 333.78662, 333.82156, 333.85406, 333.88364, 333.90976, 333.932, 333.9501, 333.96402, 333.97388, 333.9797, 333.98178, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 335.4393, 335.4684, 335.49155, 335.50797, 335.5169, 335.51758, 335.51004, 335.49564, 335.476, 335.4528, 335.42725, 335.40033, 335.37286, 335.3456, 335.3193, 335.29434, 335.2711, 335.24997, 335.2312, 335.21487, 335.201, 335.18958, 335.1806, 335.17395, 335.1695, 335.1671, 335.1667, 335.168, 335.17084, 335.17505, 335.1804, 335.18655, 335.1933, 335.20032, 335.20737, 335.2142, 335.2206, 335.22644, 335.23148, 335.23547, 335.2383, 335.23975, 335.2399, 335.23907, 335.23688, 335.2333, 335.22845, 335.22247, 335.21555, 335.2078, 335.19943, 335.19058, 335.1813, 335.17175, 335.16196, 335.15204, 335.14206, 335.132, 335.12192, 335.11182, 335.10162, 335.09125, 335.08066, 335.0753, 335.06448, 335.05365, 335.04294, 335.03244, 335.02237, 335.01297, 335.0044, 334.99683, 334.99042, 334.9852, 334.9813, 334.97876, 334.97757, 334.97766, 334.97897, 334.98145, 334.9849, 334.98917, 334.9941, 334.99954, 335.00543, 335.01172, 335.01834, 335.0253, 335.0326, 335.04025, 335.04828, 335.0567, 335.06558, 335.07587, 335.08575, 335.0961, 335.10687, 335.11795, 335.12927, 335.14078, 335.15234, 335.16388, 335.1753, 335.18652, 335.1976, 335.20856, 335.2194, 335.23013, 335.24078, 335.2513, 335.2617, 335.2719, 335.28198, 335.29196, 335.3018, 335.30667, 335.3163, 335.3258, 335.33517, 335.34436, 335.3533, 335.362, 335.37042, 335.37845, 335.3861, 335.39334, 335.40015, 335.4065, 335.4124, 335.41794, 335.42313, 335.42798, 335.4326, 335.43698, 335.4412, 335.4453, 335.44934, 335.45334, 335.45737, -999.0, -999.0, 335.47046, 335.47568, 335.48157, 335.48825, 335.4958, 335.5042, 335.5088, 335.51868, 335.52942, -999.0, -999.0, -999.0, -999.0, -999.0, 335.60516, 335.6116, 335.62405, 335.63574, 335.64627, 335.65536, 335.66284, 335.6686, 335.67255, 335.67462, 335.67477, 335.6731, 335.6716, 335.66727, 335.66122, 335.65344, 335.64395, 335.6327, 335.61978, 335.60556, 335.5904, 335.57474, 335.55902, 335.5513, 335.53656, 335.52322, 335.5119, 335.5033, 335.49826, 335.49756, 335.50204, 335.51205, -999.0, 335.55154, 335.5792, 335.61148, 335.6468, 335.68347, 335.7199, 335.75525, 335.7891, 335.82098, 335.85052, 335.8776, 335.8902, 335.91354, 335.93442, 335.95288, 335.96924, 335.98376, 335.99683, 336.00864, 336.0194, 336.02927, 336.0384, 336.0427, 336.0508, 336.05823, 336.06482, 336.0706, 336.07544, 336.07935, 336.0823, 336.0843, 336.0853, 336.08536, 336.08502, 336.0837, 336.08148, 336.0784, 336.0744, 336.06952, 336.06378, 336.0572, 336.04974, 336.04147, 336.03702, 336.0274, 336.0168, 336.0051, 335.9922, 335.97818, 335.96323, 335.94754, 335.93137, 335.91498, 335.8988, 335.8832, 335.86865, 335.8559, 335.84598, 335.83997, 335.8389, 335.84314, 335.85266, 335.86746, 335.88742, 335.89917, 335.92538, 335.95428, 335.9847, 336.01566, 336.04678, 336.07788, 336.1087, 336.13904, 336.16882, 336.19803, 336.22665, 336.25467, 336.2822, 336.3094, 336.3364, 336.36334, 336.39026, 336.41718, 336.44412, 336.47107, 336.49792, 336.52457, 336.55087, 336.57666, 336.60184, 336.62616, 336.64948, 336.67163, 336.69232, 336.71136, 336.7202, 336.73633, 336.75034, 336.76224, 336.772, 336.77972, 336.7854, 336.78928, 336.79147, 336.79218, 336.79202, 336.7908, 336.78857, 336.78552, 336.78183, 336.77762, 336.77307, 336.7683, 336.76346, 336.7587, 336.75372, 336.74954, 336.74588, 336.74292, 336.7408, 336.73975, 336.73987, 336.7413, 336.7441, 336.74838, 336.7542, 336.75772, 336.76587, 336.77557, 336.78683, 336.79956, 336.81372, 336.82922, 336.84598, 336.86392, 336.88293, 336.90295, 336.9133, 336.93466, 336.957, 336.98038, 337.00488, 337.0307, 337.05792, 337.0868, 337.11746, 337.15012, 337.18478, 337.20288, 337.24063, 337.2805, 337.3223, 337.36578, 337.41064, 337.45667, 337.5034, 337.55038, 337.59714, 337.64325, 337.66592, 337.71042, 337.75354, 337.79504, 337.83475, 337.87268, 337.90884, 337.94333, 337.97617, 338.00735, 338.03693, 338.05112, 338.07834, 338.10394, 338.12784, 338.14993, 338.17014, 338.18835, 338.20444, 338.21823, 338.2296, 338.23853, 338.24496, 338.24887, 338.2503, 338.24933, 338.24615, 338.24094, 338.23392, 338.22537, 338.21555, 338.2048, 338.19345, 338.18185, 338.17047, 338.15976, 338.1502, 338.1422, 338.13626, 338.13272, 338.13208, 338.13452, 338.1369, 338.14398, 338.15414, 338.16733, 338.1833, 338.20166, 338.22214, 338.24432, 338.2679, 338.29498, 338.32028, 338.34583, 338.37137, 338.39667, 338.42148, 338.44553, 338.46884, 338.49136, 338.5131, 338.534, 338.54413, 338.5638, 338.58273, 338.60086, 338.61826, 338.6349, 338.65082, 338.66605, 338.68057, 338.69437, 338.7074, 338.71964, 338.73105, 338.74155, 338.75104, 338.75946, 338.7668, 338.77325, 338.77887, 338.78372, 338.78802, 338.78998, 338.7937, 338.7972, 338.8007, 338.8043, 338.8082, 338.81253, 338.81744, 338.82303, 338.8293, 338.83276, 338.84024, 338.84854, 338.85773, 338.86777, 338.8787, 338.89056, 338.90338, 338.91718, 338.932, 338.94778, 338.96442, 338.97302, -999.0, 339.00888, 339.02744, 339.04617, 339.065, 339.0837, 339.10226, 339.12054, 339.13852, 339.1561, 339.17325, 339.18994, 339.20612, 339.2218, 339.237, 339.2519, 339.2665, 339.28098, 339.2954, 339.30264, 339.31723, 339.33203, 339.34717, 339.36255, 339.37823, 339.39413, 339.41022, 339.42624, 339.44205, -999.0, 339.4723, 339.47952, 339.4937, 339.50748, 339.5209, 339.534, 339.54684, 339.55948, 339.572, 339.5843, 339.59637, 339.60815, 339.6196, 339.63068, -999.0, -999.0, -999.0, -999.0, 339.67786, 339.68552, 339.6926, 339.69656, 339.70282, 339.70862, 339.714, 339.71896, 339.72342, 339.7272, 339.7303, 339.73248, 339.73367, 339.73383, 339.73312, 339.73102, 339.72745, 339.72235, 339.71573, 339.70755, 339.69794, 339.687, 339.6749, 339.6617, 339.64758, 339.6326, 339.61685, 339.60052, -999.0, -999.0, -999.0, -999.0, -999.0, 339.50906, 339.50107, 339.48544, 339.47046, -999.0, -999.0, -999.0, 339.42, 339.41043, -999.0, -999.0, 339.3911, 339.38846, 339.38815, 339.39047, 339.39597, 339.40543, 339.41962, 339.4393, -999.0, 339.49426, 339.52786, 339.56448, 339.60333, 339.6438, 339.68515, 339.72678, 339.76828, 339.80948, 339.85025, 339.89047, 339.93008, 339.96924, 340.008, 340.02728, 340.06564, 340.10385, 340.14194, 340.18002}
lat =
  {39.379, -999.0, -999.0, -999.0, -999.0, -999.0, 39.37947, 39.379604, 39.379745, 39.379887, 39.380028, 39.380177, 39.38032, 39.380474, 39.380627, 39.38078, 39.380936, 39.381096, 39.381252, 39.381413, 39.381573, 39.38173, 39.38189, 39.382046, 39.382206, 39.382362, 39.38252, 39.38267, 39.382824, 39.382977, 39.38313, 39.38328, 39.383434, 39.383583, 39.383736, 39.383884, 39.384037, 39.384186, 39.38434, 39.384487, 39.38464, 39.384792, 39.38494, 39.385094, 39.385242, 39.38539, 39.38554, 39.38569, 39.385838, 39.385983, 39.386127, 39.38627, 39.386414, 39.386555, 39.386696, 39.386837, 39.38698, 39.387115, 39.387257, 39.387398, 39.387554, 39.387695, 39.387836, 39.38798, 39.388126, 39.388268, 39.388412, 39.388554, 39.3887, 39.38884, 39.388985, 39.389126, 39.38927, 39.389412, 39.389553, 39.38969, 39.389824, 39.389954, 39.390076, 39.390194, 39.390305, 39.39041, 39.39051, 39.390606, 39.390694, 39.390774, 39.390846, 39.39091, 39.390972, 39.391026, 39.39107, 39.391117, -999.0, -999.0, -999.0, -999.0, -999.0, 39.391365, 39.391407, 39.391445, 39.39149, 39.391537, 39.391586, 39.39164, 39.391693, 39.391754, 39.391815, 39.391876, 39.39194, 39.39201, 39.39208, 39.392143, 39.392212, 39.392277, 39.392345, 39.39241, 39.39247, 39.392532, 39.392593, 39.392654, 39.39271, 39.39277, 39.39283, 39.392887, 39.39295, 39.39301, 39.393074, 39.393143, 39.39321, 39.393288, 39.393368, 39.393448, 39.393536, 39.39363, 39.393726, 39.393826, 39.393932, 39.39404, 39.39415, 39.39426, 39.394375, 39.39449, 39.394608, 39.394722, 39.394836, 39.394955, 39.39507, 39.395184, 39.395298, 39.395412, 39.395523, 39.395638, 39.39575, 39.39586, 39.39597, 39.39608, 39.39619, 39.3963, 39.39641, 39.396534, 39.396645, 39.39675, 39.396862, 39.396973, 39.397083, 39.39719, 39.397297, 39.397404, 39.397507, 39.39761, 39.39771, 39.397808, 39.397903, 39.398, 39.39809, 39.398182, 39.398266, 39.398354, 39.398438, 39.398518, 39.398598, 39.398678, 39.398754, 39.398834, 39.39891, 39.39899, 39.399067, 39.399147, 39.399227, 39.399307, 39.39939, 39.399475, 39.39956, 39.399647, 39.399734, 39.399826, 39.39992, 39.400017, 39.400112, 39.400215, 39.40032, 39.40042, 39.400528, 39.40064, 39.400753, 39.400867, 39.40098, 39.4011, 39.401222, 39.401344, 39.401466, 39.40159, 39.40171, 39.40183, 39.40195, 39.40207, 39.402184, 39.402298, 39.40241, 39.40252, 39.402622, 39.402725, 39.402824, 39.40292, 39.40301, 39.403103, 39.403187, 39.403275, 39.403355, 39.40344, 39.40352, 39.4036, 39.403675, 39.403755, 39.403835, 39.40391, 39.403996, 39.404076, 39.404156, 39.40424, 39.404324, 39.404408, 39.404495, 39.404583, 39.40467, 39.40476, 39.40485, 39.40494, 39.40503, 39.40512, 39.405212, 39.4053, 39.40539, 39.40548, 39.405567, 39.405655, 39.405743, 39.405827, 39.40591, 39.40599, 39.40607, 39.40615, 39.406227, 39.40631, 39.406384, 39.406456, 39.406525, 39.406593, 39.40666, 39.406727, 39.40679, 39.406857, 39.406918, 39.406982, 39.407047, 39.40711, 39.407173, 39.407238, 39.407303, 39.407368, 39.407433, 39.407497, 39.407566, 39.40763, 39.4077, 39.407764, 39.40783, 39.407898, 39.407963, 39.408028, 39.408092, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 39.41282, 39.412895, 39.412975, 39.413055, 39.413143, 39.41323, 39.41332, 39.413418, 39.41351, 39.4136, 39.41369, 39.41378, 39.413868, 39.413956, 39.414043, 39.414127, 39.41421, 39.41429, 39.41437, 39.414448, 39.414528, 39.414604, 39.41468, 39.414757, 39.414833, 39.41491, 39.41499, 39.415073, 39.415157, 39.415245, 39.415333, 39.41543, 39.415524, 39.415623, 39.415726, 39.41583, 39.415936, 39.416046, 39.416157, 39.41627, 39.41638, 39.416496, 39.41661, 39.416725, 39.416836, 39.416946, 39.417057, 39.417164, 39.41727, 39.417377, 39.41748, 39.41758, 39.41768, 39.417774, 39.41787, 39.417965, 39.418056, 39.418144, 39.418236, 39.418324, 39.41841, 39.418495, 39.418583, 39.418667, 39.418755, 39.41884, 39.418922, 39.419003, 39.419086, 39.419167, 39.41925, 39.41933, 39.419407, 39.419483, 39.41956, 39.419632, 39.4197, 39.41977, 39.419834, 39.4199, 39.419956, 39.420013, 39.420063, 39.420113, 39.42016, 39.4202, 39.42024, 39.420277, 39.42031, 39.42034, 39.420372, 39.4204, 39.420425, 39.420452, 39.42048, 39.4205, 39.42053, 39.42055, 39.420578, 39.420605, 39.42063, 39.42066, 39.420685, 39.42071, 39.42074, 39.420765, 39.42079, 39.42082, 39.420845, 39.42087, 39.4209, 39.420925, 39.42095, 39.420975, 39.421, 39.421024, 39.421047, 39.421066, 39.421085, 39.421104, 39.42112, 39.421135, 39.421146, 39.421158, 39.421165, 39.42117, 39.42117, 39.42117, 39.42117, 39.42116, 39.421158, 39.42115, 39.421143, 39.42113, 39.421124, 39.421116, 39.421104, 39.421097, 39.421093, 39.421085, 39.421085, 39.42108, 39.42108, 39.42108, 39.421085, 39.42109, 39.421093, 39.4211, 39.421104, 39.421112, 39.42112, 39.42113, 39.42114, 39.421146, 39.421158, 39.421165, 39.421177, 39.42119, 39.421196, 39.421207, 39.421223, 39.421234, 39.42125, 39.421265, 39.42128, 39.4213, 39.421318, 39.421337, 39.421356, 39.42138, 39.421402, 39.421425, 39.421448, 39.421467, 39.42149, 39.421505, 39.421524, 39.42154, 39.42155, 39.42156, 39.421566, 39.42157, 39.42157, 39.421566, 39.42156, 39.42155, 39.42154, 39.421528, 39.421513, 39.421497, 39.42148, 39.42146, 39.42144, 39.42142, 39.421402, 39.42138, 39.421356, 39.42133, 39.421303, 39.421276, 39.42124, 39.421207, 39.421165, 39.421124, 39.421074, 39.42102, 39.42096, 39.4209, 39.42083, 39.420753, 39.420677, 39.420586, 39.4205, 39.420414, 39.420322, 39.42023, 39.420135, 39.42004, 39.419945, 39.41985, 39.419758, 39.419662, 39.419575, -999.0, -999.0, -999.0, 39.41923, 39.41915, 39.41907, 39.418995, 39.418922, 39.418846, 39.418774, 39.4187, 39.41863, 39.418556, 39.41848, 39.418404, 39.418324, 39.418243, 39.41816, 39.41807, 39.417984, 39.41789, 39.417793, 39.417694, 39.41759, 39.41749, 39.41738, 39.41727, 39.41716, 39.417046, 39.416927, 39.416813, 39.416695, 39.416576, 39.41646, 39.41634, 39.416225, 39.416107, 39.415993, 39.41588, 39.415768, 39.415653, 39.415546, 39.415436, 39.41533, 39.415222, 39.415115, 39.41501, 39.4149, 39.4148, 39.414692, 39.414585, 39.41448, 39.41437, 39.41426, 39.414154, 39.414043, 39.413933, 39.413822, 39.413715, 39.413605, 39.413494, 39.413383, 39.413273, 39.413162, 39.41305, 39.41294, 39.41283, 39.412716, 39.4126, 39.412483, 39.41236, 39.41224, 39.412113, 39.411983, 39.41185, 39.411713, 39.41157, 39.411427, 39.411278, 39.411125, 39.410957, 39.410797, 39.41064, 39.41048, 39.41032, 39.41016, 39.409996, 39.40984, 39.40968, 39.409523, 39.40937, 39.409218, 39.40907, 39.408924, 39.408783, 39.40864, 39.408504, 39.40837, 39.40824, 39.40811, 39.407986, 39.407864, 39.407745, 39.407627, 39.407513, 39.407402, 39.40729, 39.40718, 39.407078, 39.406975, 39.40687, 39.40677, 39.40667, 39.40657, 39.40647, 39.406372, 39.406273, 39.406174, 39.40607, 39.405968, 39.40586, 39.405754, 39.405643, 39.405533, 39.40542, 39.4053, 39.40518, 39.405064, 39.40494, 39.404816, 39.404694, 39.404568, 39.40444, 39.404312, 39.404182, 39.404053, 39.403923, 39.40379, 39.403656, 39.403522, 39.403385, 39.403244, 39.403103, 39.40296, 39.402813, 39.402664, 39.40251, 39.402355, 39.4022, 39.40204, 39.401875, 39.40171, 39.401543, 39.40137, 39.401203, 39.40103, 39.40086, 39.40069, 39.400517, 39.400345, 39.400173, 39.4, 39.399834, 39.399666, 39.3995, 39.399338, 39.399174, 39.39901, 39.39885, 39.39869, 39.39853, 39.39837, 39.398212, 39.398052, 39.397896, 39.39774, 39.397583, 39.397427, 39.397274, 39.397118, 39.396965, 39.39681, 39.39664, 39.39649, 39.396336, 39.396183, 39.39603, 39.395878, 39.39572, 39.39557, 39.395416, 39.395264, 39.39511, 39.394955, 39.394802, 39.394646, 39.39449, 39.394333, 39.394176, 39.39402, 39.393864, 39.393707, 39.393547, 39.39339, 39.393234, 39.393078, 39.39292, 39.39276, 39.392605, 39.39245, 39.392292, 39.392136, 39.39198, 39.391823, 39.391666, 39.391506, 39.391346, 39.391186, 39.391026, 39.390858, 39.390694, 39.390526, 39.390354, 39.390182, 39.390007, 39.38983, 39.389652, 39.389473, 39.389294, 39.389114, 39.38894, 39.38876, 39.388584, 39.38841, 39.388325, 39.388153, 39.38799, 39.387825, 39.38767, 39.387512, 39.387356, 39.387207, 39.38706, 39.386913, 39.38677, 39.386623, 39.38648, 39.386337, 39.386192, 39.386047, 39.3859, 39.385754, 39.385605, 39.385452, 39.3853, 39.385147, 39.38499, 39.38484, 39.38468, 39.384525, 39.384365, 39.38421, 39.384052, 39.3839, 39.383743, 39.383587, 39.383434, 39.38328, 39.38313, 39.38298, 39.382828, 39.38268, 39.382526, 39.382378, 39.38223, 39.382076, 39.381924, 39.38177, 39.38162, 39.381466, 39.38131, 39.38115, 39.380993, 39.380833, 39.380657, 39.380493, 39.38033, 39.380165, 39.38, 39.379837, 39.379673, 39.37951, 39.379345, 39.37918, 39.379017, 39.378857, 39.378693, 39.378532, 39.378372, 39.37821, 39.37805, 39.37789, 39.37773, 39.37757, 39.377415, 39.377254, 39.377098, 39.376938, 39.37678, 39.37662, 39.37646, 39.376305, 39.376144, 39.375984, 39.375828, 39.375668, 39.37551, 39.37535, 39.375195, 39.375034, 39.374878, 39.37472, 39.374565, 39.37441, 39.374252, 39.374096, 39.373943, 39.373787, 39.373627, 39.37347, 39.373314, 39.373154, 39.372993, 39.37283, 39.372665, 39.372498, 39.37233, 39.37216, 39.37199, 39.371815, 39.37164, 39.371464, 39.37129, 39.37111, 39.37093, 39.37075, 39.370575, 39.370396, 39.370216, 39.37004, 39.36986, 39.36969, 39.369514, 39.369343, 39.369175, 39.369007, 39.36884, 39.368675, 39.368507, 39.368347, 39.368183, 39.368023, 39.36786, 39.3677, 39.36754, 39.367374, 39.367214, 39.367054, 39.36689, 39.36673, 39.366566, 39.3664, 39.36624, 39.366077, 39.365913, 39.365753, 39.36559, 39.365425, 39.365265, 39.365105, 39.36494, 39.36478, 39.36462, 39.364456, 39.364292, 39.364132, 39.36395, 39.363785, 39.363617, 39.36345, 39.36328, 39.36311, 39.362934, 39.36276, 39.362583, 39.362404, 39.36222, 39.36204, 39.36186, 39.36167, 39.36149, 39.3613, 39.36112, 39.36093, 39.360744, 39.36056, 39.360374, 39.36019, 39.36001, 39.359825, 39.359642, 39.359463, 39.35928, 39.359097, 39.358917, 39.358738, 39.358555, 39.358376, 39.358192, 39.358013, 39.35783, 39.35765, 39.357468, 39.357285, 39.357105, 39.356922, 39.35674, 39.356647, 39.356464, 39.35628, 39.3561, 39.355915, 39.355736, 39.355553, 39.355373, 39.355194, 39.35502, 39.35484, 39.354664, 39.35449, 39.354313, 39.35414, 39.35397, 39.353798, 39.353626, 39.353455, 39.353287, 39.353115, 39.352943, 39.35277, 39.3526, 39.35243, 39.352253, 39.352077, 39.3519, 39.351723, 39.35154, 39.35136, 39.351177, 39.350994, 39.35081, 39.350624, 39.35044, 39.350254, 39.350067, 39.349884, 39.3497, 39.349514, 39.34933, 39.34915, 39.34897, 39.34879, 39.34861, 39.34843, 39.348255, 39.348076, 39.3479, 39.34773, 39.347553, 39.347378, 39.347206, 39.34703, 39.34686, 39.346687, 39.34651, 39.34634, 39.346165, 39.34599, 39.345814, 39.34564, 39.345463, 39.345284, 39.345104, 39.34492, 39.344738, 39.344555, 39.344368, 39.34418, 39.343994, 39.343784, 39.343594, 39.343403, 39.34321, 39.343018, 39.342823, 39.34263, 39.342438, 39.342243, 39.342052, 39.34186, 39.34167, 39.34148, 39.341293, 39.341106, 39.34092, 39.340733, 39.34055, 39.340366, 39.340187, 39.340004, 39.339916, 39.339737, 39.339558, 39.33938, 39.3392, 39.339024, 39.338844, 39.33867, 39.33849, 39.33831, 39.338135, 39.337955, 39.33778, 39.3376, 39.33742, 39.337242, 39.337063, 39.336884, 39.336704, 39.33652, 39.33634, 39.33616, 39.335976, 39.335793, 39.335613, 39.33543, 39.335247, 39.335068, 39.33489, 39.33471, 39.33453, 39.334354, 39.334183, 39.33401, 39.33384, 39.33367, 39.333508, 39.333344, 39.33318, 39.33302, 39.33286, 39.332703, 39.332542, 39.332386, 39.33223, 39.332073, 39.331917, 39.33176, 39.3316, 39.331444, 39.331284, 39.331123, 39.33096, 39.3308, 39.330635, 39.330467, 39.330303, 39.330135, 39.329967, 39.3298, 39.32963, 39.329464, 39.329296, 39.32913, 39.32896, 39.328793, 39.328625, 39.32846, 39.328293, 39.32813, 39.327965, 39.3278, 39.327637, 39.32747, 39.327305, 39.32714, 39.326977, 39.326813, 39.32665, 39.326485, 39.326317, 39.326153, 39.32605, 39.325882, 39.325714, 39.325546, 39.325375, 39.325207, 39.325035, 39.324863, 39.324688, 39.324516, 39.32434, 39.324165, 39.32399, 39.323814, 39.323635, 39.32346, 39.323284, 39.323105, 39.32293, 39.322754, 39.322575, 39.3224, 39.322224, 39.32205, 39.321873, 39.3217, 39.321526, 39.321354, 39.32118, 39.321007, 39.320835, 39.320663, 39.32049, 39.320316, 39.320145, 39.319973, 39.3198, 39.31963, 39.319458, 39.319283, 39.31911, 39.318935, 39.31876, 39.318584, 39.31841, 39.31823, 39.318054, 39.317875, 39.317696, 39.317516, 39.317337, 39.317158, 39.316975, 39.316795, 39.316612, 39.31643, 39.316246, 39.316067, 39.315884, 39.3157, 39.315517, 39.31534, 39.315155, 39.314972, 39.314793, 39.31461, 39.314426, 39.314247, 39.314064, 39.31388, 39.3137, 39.31352, 39.313335, 39.313152, 39.312973, 39.31279, 39.312607, 39.312424, 39.31224, 39.312057, 39.311874, 39.31169, 39.3116, 39.311417, 39.311234, 39.311054, 39.31087, 39.31069, 39.31051, 39.31033, 39.31015, 39.30997, 39.309772, 39.309593, 39.309414, 39.309235, 39.309055, 39.308876, 39.308697, 39.308517, 39.30834, 39.30816, 39.30798, 39.3078, 39.30762, 39.30744, 39.307262, 39.307083, 39.306904, 39.306725, 39.30655, 39.306374, 39.306194, 39.30602, 39.305843, 39.305668, 39.305492, 39.305317, 39.30514, 39.304966, 39.30479, 39.30461, 39.304432, 39.304253, 39.30407, 39.303886, 39.303703, 39.303516, 39.30333, 39.303143, 39.302956, 39.30277, 39.302578, 39.302387, 39.3022, 39.30201, 39.30182, 39.301632, 39.30144, 39.301254, 39.301067, 39.30088, 39.300697, 39.300602, 39.30042, 39.300236, 39.300053, 39.29987, 39.299686, 39.299507, 39.299324, 39.29914, 39.29896, 39.29878, 39.298595, 39.298416, 39.298233, 39.298054, 39.29787, 39.29769, 39.29751, 39.29733, 39.29715, 39.29697, 39.29679, 39.296616, 39.296436, 39.29626, 39.296085, 39.29591, 39.295734, 39.295563, 39.29539, 39.29522, 39.295048, 39.294876, 39.29471, 39.29454, 39.294376, 39.29421, 39.294044, 39.29388, 39.29372, 39.29356, 39.2934, 39.293324, 39.293167, 39.29301, 39.29286, 39.292706, 39.292557, 39.292408, 39.29226, 39.292114, 39.29197, 39.29181, 39.291664, 39.291523, 39.291378, 39.291237, 39.291096, 39.290955, 39.290813, 39.290676, 39.290535, 39.290398, 39.29026, 39.290123, 39.289986, 39.28985, 39.289715, 39.28958, 39.289448, 39.289314, 39.28918, 39.28905, 39.28892, 39.28879, 39.288666, 39.288536, 39.28841, 39.28829, 39.288162, 39.28804, 39.28792, 39.287804, 39.287685, 39.28757, 39.287457, 39.287346, 39.28724, 39.287132, 39.28703, 39.286926, 39.286827, 39.28673, 39.28664, 39.28655, 39.28646, 39.286377, 39.286293, 39.286213, 39.286133, 39.286057, 39.28598, 39.285908, 39.285835, 39.285763, 39.285694, 39.285625, 39.285557, 39.28549, 39.285423, 39.28536, 39.285294, 39.285233, 39.285168, 39.285107, 39.285046, 39.284985, 39.284924, 39.284863, 39.2848, 39.28474, 39.284676, 39.284615, 39.284554, 39.28449, 39.284428, 39.284363, 39.2843, 39.284237, 39.284176, 39.284115, 39.284054, 39.283993, 39.28393, 39.283875, 39.28382, 39.283768, 39.283714, 39.283665, 39.283615, 39.28357, 39.283527, 39.283485, 39.283443, 39.283424, 39.283386, 39.283348, 39.28331, 39.283276, 39.283237, 39.2832, 39.283165, 39.283127, 39.283085, 39.283043, 39.283, 39.282963, 39.28292, 39.28288, 39.282833, 39.28279, 39.28275, 39.282703, 39.28266, 39.282616, 39.282574, 39.28253, 39.28249, 39.282448, 39.282406, 39.282364, 39.282322, 39.282276, 39.282234, 39.282192, 39.282146, 39.2821, 39.28205, 39.282005, 39.281956, 39.281902, 39.281853, 39.2818, 39.281742, 39.28169, 39.28163, 39.281574, 39.281517, 39.281456, 39.2814, 39.281338, 39.281277, 39.281216, 39.281155, 39.281094, 39.281033, 39.28097, 39.28091, 39.28085, 39.28079, 39.280727, 39.280666, 39.280605, 39.280544, 39.28048, 39.28042, 39.280357, 39.280296, 39.280235, 39.280174, 39.280113, 39.280052, 39.27999, 39.27993, 39.27987, 39.279808, 39.279747, 39.279686, 39.279625, 39.279564, 39.279503, 39.279446, 39.27939, 39.27933, 39.279274, 39.279217, 39.27919, 39.279137, 39.279087, 39.279034, 39.278984, 39.278934, 39.27889, 39.27884, 39.278793, 39.278748, 39.2787, 39.278656, 39.27861, 39.278564, 39.27852, 39.278473, 39.278427, 39.27838, 39.27833, 39.278286, 39.278236, 39.278183, 39.278133, 39.278076, 39.278023, 39.277966, 39.277905, 39.277843, 39.27778, 39.27771, 39.27764, 39.277565, 39.277493, 39.277412, 39.27733, 39.277245, 39.277153, 39.27706, 39.276962, 39.276863, 39.27676, 39.276646, 39.27654, 39.27643, 39.276318, 39.276203, 39.27609, 39.275974, 39.27586, 39.275745, 39.27563, 39.275517, 39.275406, 39.27529, 39.275185, 39.275074, 39.274967, 39.274864, 39.27476, 39.274662, 39.274567, 39.27447, 39.27438, 39.27429, 39.274197, 39.274113, 39.274025, 39.273945, 39.27386, 39.27378, 39.2737, 39.273624, 39.27355, 39.27347, 39.273396, 39.27332, 39.273243, 39.27317, 39.273094, 39.273018, 39.27294, 39.272865, 39.27279, 39.27271, 39.272633, 39.272552, 39.272472, 39.272392, 39.27231, 39.27223, 39.272144, 39.272064, 39.27198, 39.271896, 39.271816, 39.271732, 39.27165, 39.271564, 39.27148, 39.271397, 39.271313, 39.27123, 39.271145, 39.27106, 39.270973, 39.270885, 39.270798, 39.27071, 39.270622, 39.27053, 39.270443, 39.27035, 39.27026, 39.27017, 39.270073, 39.26998, 39.269886, 39.26979, 39.269695, 39.2696, 39.2695, 39.2694, 39.269302, 39.2692, 39.269096, 39.268993, 39.268887, 39.26878, 39.26867, 39.268555, 39.26844, 39.268322, 39.268204, 39.26808, 39.267956, 39.267826, 39.267693, 39.26756, 39.26742, 39.267284, 39.267143, 39.267, 39.266857, 39.266697, 39.266556, 39.26641, 39.26627, 39.26613, 39.26599, 39.265858, 39.265724, 39.265594, 39.26547, 39.265347, 39.265224, 39.265106, 39.264988, 39.26487, 39.26475, 39.264637, 39.26452, 39.264397, 39.26428, 39.264153, 39.264027, 39.2639, 39.263767, 39.263634, 39.2635, 39.26336, 39.26322, 39.26308, 39.26294, 39.2628, 39.262657, 39.262516, 39.26238, 39.26224, 39.262108, 39.261974, 39.261845, 39.26172, 39.261593, 39.26147, 39.26135, 39.26123, 39.261116, 39.261, 39.260887, 39.26078, 39.26067, 39.260567, 39.26046, 39.26036, 39.26026, 39.260166, 39.260075, 39.259987, 39.2599, 39.259815, 39.25973, 39.259655, 39.259575, 39.2595, 39.259422, 39.25935, 39.259274, 39.259197, 39.259117, 39.259037, 39.258957, 39.25887, 39.25878, 39.25869, 39.258595, 39.258495, 39.258446, 39.258343, 39.258236, 39.258125, 39.25802, 39.257904, 39.257793, 39.257683, 39.257572, 39.257465, 39.257412, 39.257305, 39.257206, 39.257107, 39.257008, 39.256916, 39.25682, 39.256733, 39.25664, 39.25655, 39.25645, 39.25636, 39.256268, 39.25617, 39.25607, 39.255966, 39.25586, 39.25575, 39.255634, 39.255516, 39.255394, 39.255272, 39.25515, 39.255028, 39.2549, 39.25478, 39.25466, 39.254547, 39.254433, 39.254326, 39.254272, 39.25417, 39.254074, 39.25398, 39.25389, 39.2538, 39.253716, 39.253628, 39.253544, 39.253456, 39.253372, 39.253326, 39.25324, 39.253147, 39.25305, 39.252953, 39.252853, 39.25275, 39.252644, 39.252533, 39.252422, 39.252304, 39.252247, 39.25213, 39.25201, 39.251892, 39.251774, 39.251656, 39.251537, 39.251423, 39.251312, 39.2512, 39.251095, 39.25099, 39.250893, 39.250793, 39.2507, 39.25061, 39.250523, 39.250435, 39.25035, 39.25027, 39.250187, 39.250107, 39.250027, 39.249943, 39.24986, 39.249775, 39.249687, 39.249596, 39.2495, 39.249405, 39.249306, 39.249207, 39.2491, 39.248993, 39.248886, 39.248775, 39.24866, 39.248547, 39.248436, 39.24832, 39.248207, 39.248096, 39.24804, 39.24793, 39.24782, 39.247715, 39.24761, 39.247505, 39.247406, 39.247307, 39.247208, 39.247112, 39.247063, 39.246967, 39.24687, 39.246773, 39.246677, 39.24658, 39.24648, 39.246376, 39.246273, 39.246166, 39.24606, 39.246006, 39.245895, 39.245785, 39.245674, 39.245564, 39.24545, 39.24534, 39.245228, 39.245117, 39.245064, 39.244953, 39.244892, 39.244785, 39.244686, 39.244583, 39.244488, 39.244392, 39.244297, 39.2442, 39.24411, 39.244022, 39.24393, 39.243843, 39.24375, 39.243664, 39.243576, 39.243484, 39.243397, 39.243305, 39.243214, 39.243122, 39.243027, 39.24293, 39.24284, 39.242744, 39.242645, 39.24255, 39.24245, 39.24235, 39.242252, 39.242153, 39.242054, 39.242004, 39.2419, 39.2418, 39.241695, 39.241592, 39.24149, 39.241386, 39.24128, 39.241173, 39.241066, 39.24096, 39.240852, 39.240746, 39.240635, 39.240524, 39.240414, 39.240307, 39.240196, 39.240086, 39.239975, 39.23987, 39.239758, 39.23965, 39.23954, 39.239433, 39.239323, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 39.219875, 39.219738, 39.2196, 39.21946, 39.21932, 39.21918, 39.21904, 39.2189, 39.218758, 39.21862, 39.21848, 39.21834, 39.2182, 39.218063, 39.21793, 39.217793, 39.217655, 39.21752, 39.21739, 39.217255, 39.217117, 39.216984, 39.21685, 39.216713, 39.21658, 39.216442, 39.216305, 39.216167, 39.21603, 39.215893, 39.21575, 39.21561, 39.215473, 39.215332, 39.21519, 39.21505, 39.21491, 39.214764, 39.214622, 39.21448, 39.214336, 39.214195, 39.214127, 39.213985, 39.213844, 39.213703, 39.213562, 39.213425, 39.213287, 39.21315, 39.213013, 39.212875, 39.212738, 39.212605, 39.21247, 39.212334, 39.2122, 39.212067, 39.21193, 39.211796, 39.21166, 39.211525, 39.211388, 39.21132, 39.21118, 39.211044, 39.210903, 39.210766, 39.21063, 39.210487, 39.21035, 39.210213, 39.21007, 39.209934, 39.209797, 39.20966, 39.209522, 39.209385, 39.209244, 39.209106, 39.20897, 39.20883, 39.208694, 39.208557, 39.20842, 39.208282, 39.20814, 39.208004, 39.207863, 39.20772, 39.20758, 39.207436, 39.207294, 39.207138, 39.206993, 39.20685, 39.206707, 39.206562, 39.206417, 39.206276, 39.206135, 39.205994, 39.205856, 39.20572, 39.20558, 39.20545, 39.20532, 39.205185, 39.20506, 39.204933, 39.20481, 39.20469, 39.204567, 39.204453, 39.204334, 39.204277, 39.204163, 39.20405, 39.203938, 39.203823, 39.203712, 39.203598, 39.203487, 39.203373, 39.20326, 39.203144, 39.203026, 39.202908, 39.20279, 39.202667, 39.20254, 39.20242, 39.20229, 39.20216, 39.20203, 39.201897, 39.201763, 39.20163, 39.201492, 39.201355, 39.201214, 39.201077, 39.200935, 39.200794, 39.200653, 39.20051, 39.200363, 39.20029, 39.200146, 39.199997, 39.19985, 39.199696, 39.199543, 39.19939, 39.199234, 39.199074, 39.198997, 39.198837, 39.198673, 39.19851, 39.19835, 39.198185, 39.19802, 39.197853, 39.19769, 39.197525, 39.19736, 39.19728, 39.197117, 39.196957, 39.196793, 39.196632, 39.196472, 39.196312, 39.196156, 39.195995, 39.19584, 39.195683, 39.195602, 39.19545, 39.195293, 39.19514, 39.19499, 39.194836, 39.194683, 39.194534, 39.194386, 39.19422, 39.194073, 39.193928, 39.19378, 39.193634, 39.19349, 39.193344, 39.193195, 39.19305, 39.192905, 39.19276, 39.19261, 39.19254, 39.19239, 39.192238, 39.19209, 39.191933, 39.19178, 39.191624, 39.191463, 39.191303, 39.191143, 39.19098, 39.1909, 39.19073, 39.190567, 39.190403, 39.190235, 39.19007, 39.189903, 39.18974, 39.18958, 39.18942, 39.18926, 39.189182, 39.189026, 39.188877, 39.188725, 39.18858, 39.188435, 39.188293, 39.188152, 39.188015, 39.18788, 39.187813, 39.187683, 39.18755, 39.18742, 39.187286, 39.187157, 39.187023, 39.18689, 39.186756, 39.186623, 39.186485, 39.186344, 39.186207, 39.18606, 39.18592, 39.185776, 39.18563, 39.185486, 39.185337, 39.185192, 39.185047, 39.184975, 39.184834, 39.18469, 39.184547, 39.184406, 39.184265, 39.184124, 39.183987, 39.183846, 39.183704, 39.183563, 39.18342, 39.183273, 39.18313, 39.18298, 39.182827, 39.18268, 39.18252, 39.18237, 39.182213, 39.182056, 39.1819, 39.18174, 39.181583, 39.181427, 39.18127, 39.181114, 39.18096, 39.18081, 39.18066, 39.18051, 39.18044, 39.180298, 39.180157, 39.18002, 39.179882, 39.179745, 39.17961, 39.17948, 39.17935, 39.179222, 39.179157, 39.179028, 39.1789, 39.178772, 39.178642, 39.178513, 39.178383, 39.178253, 39.178123, 39.177994, 39.17785, 39.177715, 39.177586, 39.177456, 39.177322, 39.177197, 39.177067, 39.17694, 39.176815, 39.17669, 39.176567, 39.176506, 39.176388, 39.176266, 39.17615, 39.176033, 39.17592, 39.175804, 39.175694, 39.175583, 39.175472, 39.17536, 39.17531, 39.1752, 39.175095, 39.174988, 39.17488, 39.174778, 39.17467, 39.17457, 39.174465, 39.174362, 39.17426, 39.174206, 39.174107, 39.174004, 39.1739, 39.173798, 39.1737, 39.173595, 39.173496, 39.173397, 39.173298, 39.1732, 39.17315, 39.173054, 39.17296, 39.172863, 39.172768, 39.172672, 39.172577, 39.17248, 39.172386, 39.17229, 39.17219, 39.172146, 39.172047, 39.171944, 39.171844, 39.171738, 39.171635, 39.171528, 39.171417, 39.17131, 39.1712, 39.171085, 39.170975, 39.17086, 39.17075, 39.170635, 39.170525, 39.170414, 39.170303, 39.170193, 39.170086, 39.16998, 39.169872, 39.169765, 39.169662, 39.16956, 39.169456, 39.169357, 39.169254, 39.16915, 39.16905, 39.168945, 39.168896, 39.16879, 39.168686, 39.168575, 39.16847, 39.168358, 39.168247, 39.168133, 39.16802, 39.167892, 39.167774, 39.16766, 39.16754, 39.167423, 39.16731, 39.16719, 39.167076, 39.16696, 39.16685, 39.166737, 39.166683, 39.166573, 39.166466, 39.16636, 39.166252, 39.16615, 39.166046, 39.165943, 39.16584, 39.165737, 39.165634, 39.16553, 39.16543, 39.165325, 39.165222, 39.16512, 39.165012, 39.16491, 39.164806, 39.1647, 39.164597, 39.164547, 39.16444, 39.164337, 39.164238, 39.164135, 39.164032, 39.163933, 39.16383, 39.16373, 39.16363, 39.16358, 39.163483, 39.163383, 39.163284, 39.163185, 39.163086, 39.16299, 39.16289, 39.162792, 39.162693, 39.162594, 39.162495, 39.16245, 39.16235, 39.16225, 39.162155, 39.16206, 39.161964, 39.16187, 39.161777, 39.161682, 39.16159, 39.161503, 39.16141, 39.161324, 39.161236, 39.161148, 39.16106, 39.160976, 39.160892, 39.160805, 39.16072, 39.16068, 39.160595, 39.16051, 39.160423, 39.16034, 39.160255, 39.160168, 39.160084, 39.159996, 39.159912, 39.15983, 39.15974, 39.1597, 39.159615, 39.159527, 39.159443, 39.159355, 39.15927, 39.159187, 39.159103, 39.159016, 39.15893, 39.158848, 39.158764, 39.15868, 39.158596, 39.158512, 39.15843, 39.15834, 39.158257, 39.158173, 39.15809, 39.15804, 39.157955, 39.15787, 39.157787, 39.157707, 39.157623, 39.157543, 39.157463, 39.157383, 39.157303, 39.157265, 39.157185, 39.15711, 39.15703, 39.15695, 39.15688, 39.156803, 39.156727, 39.15665, 39.156574, 39.1565, 39.156425, 39.15635, 39.156273, 39.156197, 39.15612, 39.156044, 39.155964, 39.155884, 39.155804, 39.155724, 39.15568, 39.1556, 39.155518, 39.155434, 39.15535, 39.155266, 39.15518, 39.155098, 39.155014, 39.154926, 39.154842, 39.154755, 39.15467, 39.154587, 39.1545, 39.154415, 39.154327, 39.15424, 39.154152, 39.154064, 39.153976, 39.153893, 39.15381, 39.153732, 39.153667, 39.153618, 39.153576, 39.15355, 39.153534, 39.153526, 39.153526, 39.15353, 39.15353, 39.15353, 39.153534, 39.153534, 39.153538, -999.0}
lon =
  {-101.032, -999.0, -999.0, -999.0, -999.0, -999.0, -101.03182, -101.03178, -101.03172, -101.03167, -101.03161, -101.031555, -101.031494, -101.03143, -101.031364, -101.0313, -101.031235, -101.031166, -101.0311, -101.03102, -101.03095, -101.030876, -101.0308, -101.03072, -101.03065, -101.03057, -101.030495, -101.03042, -101.03034, -101.030266, -101.03019, -101.03011, -101.03004, -101.02997, -101.02989, -101.029816, -101.02975, -101.02967, -101.0296, -101.029526, -101.02946, -101.02939, -101.02931, -101.02924, -101.029175, -101.029106, -101.02904, -101.02897, -101.0289, -101.02883, -101.02876, -101.028694, -101.028625, -101.028564, -101.028496, -101.028435, -101.028366, -101.028305, -101.02824, -101.028175, -101.0281, -101.02804, -101.02797, -101.02791, -101.02784, -101.02778, -101.02771, -101.02764, -101.027565, -101.0275, -101.02743, -101.02735, -101.027275, -101.02721, -101.02713, -101.027054, -101.02697, -101.02689, -101.02682, -101.02674, -101.02667, -101.026596, -101.02652, -101.02645, -101.02638, -101.02631, -101.02625, -101.02619, -101.02613, -101.02607, -101.02601, -101.025955, -999.0, -999.0, -999.0, -999.0, -999.0, -101.02561, -101.02556, -101.0255, -101.02544, -101.02538, -101.02532, -101.02526, -101.0252, -101.02514, -101.02508, -101.02502, -101.024956, -101.024895, -101.02483, -101.02478, -101.02472, -101.024666, -101.02461, -101.02456, -101.024506, -101.02445, -101.0244, -101.02434, -101.024284, -101.02423, -101.02418, -101.02412, -101.024055, -101.023994, -101.02393, -101.02387, -101.0238, -101.023735, -101.02367, -101.02359, -101.02352, -101.023445, -101.02337, -101.023285, -101.02321, -101.02313, -101.02305, -101.02297, -101.02289, -101.02281, -101.022736, -101.02265, -101.02257, -101.02249, -101.02241, -101.02232, -101.02224, -101.022156, -101.022064, -101.02197, -101.02188, -101.02178, -101.02168, -101.021576, -101.02147, -101.02136, -101.02125, -101.02111, -101.02099, -101.02087, -101.02074, -101.02061, -101.02048, -101.02034, -101.0202, -101.020065, -101.01993, -101.01978, -101.019646, -101.0195, -101.019356, -101.01922, -101.01907, -101.01892, -101.018776, -101.01862, -101.01847, -101.01832, -101.01816, -101.018, -101.01783, -101.017654, -101.01748, -101.0173, -101.01712, -101.01693, -101.01674, -101.01654, -101.016335, -101.016136, -101.01592, -101.01572, -101.0155, -101.01529, -101.015076, -101.014854, -101.01464, -101.01443, -101.014206, -101.01399, -101.01377, -101.01356, -101.01334, -101.01313, -101.01292, -101.0127, -101.0125, -101.01229, -101.012085, -101.01188, -101.01167, -101.011475, -101.01128, -101.01108, -101.01088, -101.01068, -101.01048, -101.01029, -101.01009, -101.009895, -101.0097, -101.0095, -101.0093, -101.0091, -101.0089, -101.0087, -101.0085, -101.00829, -101.00809, -101.00788, -101.007675, -101.00747, -101.00726, -101.00706, -101.00685, -101.00665, -101.00645, -101.00625, -101.00605, -101.00586, -101.00567, -101.00548, -101.005295, -101.00511, -101.00493, -101.00475, -101.00458, -101.00441, -101.00424, -101.004074, -101.00391, -101.003746, -101.00358, -101.00342, -101.00326, -101.0031, -101.00294, -101.00278, -101.00262, -101.00246, -101.0023, -101.00211, -101.00195, -101.00179, -101.001625, -101.001465, -101.0013, -101.00114, -101.00097, -101.00081, -101.00065, -101.00049, -101.00033, -101.000175, -101.00002, -100.99987, -100.99972, -100.99957, -100.99943, -100.99929, -100.999146, -100.99901, -100.99887, -100.99873, -100.998604, -100.99847, -100.99834, -100.99821, -100.99807, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -100.9903, -100.990204, -100.990105, -100.990005, -100.9899, -100.989784, -100.98968, -100.98955, -100.98942, -100.989296, -100.98917, -100.98903, -100.988884, -100.98874, -100.988594, -100.98844, -100.98828, -100.98813, -100.98797, -100.98781, -100.98764, -100.98748, -100.98732, -100.98716, -100.987, -100.98684, -100.98669, -100.986534, -100.98638, -100.98624, -100.9861, -100.98596, -100.985825, -100.985695, -100.985565, -100.985435, -100.985306, -100.98518, -100.985054, -100.984924, -100.984795, -100.984665, -100.984535, -100.9844, -100.98425, -100.984116, -100.98397, -100.98382, -100.983665, -100.98351, -100.98336, -100.98321, -100.983055, -100.982895, -100.98274, -100.98259, -100.982445, -100.9823, -100.982155, -100.98202, -100.98188, -100.98174, -100.98161, -100.98148, -100.98136, -100.98124, -100.98112, -100.981, -100.98089, -100.980774, -100.98066, -100.980545, -100.98043, -100.980316, -100.9802, -100.98009, -100.97997, -100.97985, -100.97974, -100.979614, -100.97949, -100.97937, -100.97925, -100.97912, -100.97899, -100.97886, -100.97872, -100.978584, -100.97845, -100.97831, -100.978165, -100.97802, -100.977875, -100.97773, -100.977585, -100.97744, -100.977295, -100.97714, -100.977, -100.97684, -100.976685, -100.97654, -100.976395, -100.97625, -100.976105, -100.97596, -100.975815, -100.97567, -100.97553, -100.97539, -100.97525, -100.975105, -100.97497, -100.97482, -100.974686, -100.97454, -100.9744, -100.97426, -100.97411, -100.97397, -100.973816, -100.97366, -100.97351, -100.97336, -100.9732, -100.97303, -100.97287, -100.972694, -100.97253, -100.97235, -100.97217, -100.971985, -100.9718, -100.97162, -100.97143, -100.971245, -100.971054, -100.97087, -100.97069, -100.970505, -100.97032, -100.970146, -100.96997, -100.9698, -100.969635, -100.969475, -100.969315, -100.96916, -100.96901, -100.968864, -100.96872, -100.968575, -100.96843, -100.96829, -100.96815, -100.96801, -100.967865, -100.96773, -100.96758, -100.96744, -100.9673, -100.967155, -100.96701, -100.966866, -100.96673, -100.96658, -100.966446, -100.9663, -100.96616, -100.966034, -100.9659, -100.96577, -100.96564, -100.96551, -100.96538, -100.965256, -100.965126, -100.965004, -100.96488, -100.96476, -100.96463, -100.96451, -100.964386, -100.96426, -100.96413, -100.964, -100.96387, -100.96374, -100.9636, -100.96347, -100.96333, -100.963196, -100.96306, -100.96293, -100.96279, -100.96266, -100.962524, -100.962395, -100.962265, -100.962135, -100.962006, -100.96188, -100.96176, -100.96164, -100.96152, -100.961395, -100.96127, -100.96115, -100.96104, -100.960915, -100.96079, -100.960655, -100.96053, -100.9604, -100.96028, -100.96015, -100.96002, -100.95989, -100.959755, -100.959625, -100.95949, -100.95935, -100.95921, -999.0, -999.0, -999.0, -100.95866, -100.95851, -100.95837, -100.95822, -100.95808, -100.957924, -100.95778, -100.95763, -100.95747, -100.95732, -100.95717, -100.957016, -100.95687, -100.95672, -100.956566, -100.95642, -100.956276, -100.95613, -100.95599, -100.95585, -100.95571, -100.955574, -100.955444, -100.95531, -100.95517, -100.95504, -100.9549, -100.954765, -100.95462, -100.954475, -100.95433, -100.95418, -100.95402, -100.95385, -100.95368, -100.95351, -100.95333, -100.95315, -100.95296, -100.95276, -100.95256, -100.952354, -100.95215, -100.951935, -100.95172, -100.95151, -100.95129, -100.951065, -100.950836, -100.950615, -100.950386, -100.95016, -100.949936, -100.94971, -100.949486, -100.94926, -100.949036, -100.94882, -100.94861, -100.948395, -100.94819, -100.94798, -100.947784, -100.94759, -100.9474, -100.94723, -100.94705, -100.946884, -100.94672, -100.94656, -100.94641, -100.946266, -100.94613, -100.94599, -100.94586, -100.94573, -100.94561, -100.94547, -100.94535, -100.94524, -100.945114, -100.945, -100.94488, -100.944756, -100.94463, -100.94451, -100.94439, -100.94426, -100.94412, -100.943985, -100.94385, -100.9437, -100.94355, -100.943405, -100.943245, -100.94309, -100.942924, -100.942764, -100.9426, -100.94243, -100.94225, -100.94208, -100.9419, -100.94173, -100.94154, -100.94136, -100.94118, -100.94099, -100.9408, -100.940605, -100.940414, -100.940216, -100.94002, -100.93982, -100.93961, -100.9394, -100.93919, -100.93898, -100.93876, -100.93854, -100.93832, -100.93809, -100.93786, -100.93762, -100.93739, -100.93716, -100.93691, -100.936676, -100.93643, -100.93619, -100.93594, -100.93569, -100.93545, -100.9352, -100.93496, -100.934715, -100.93448, -100.93424, -100.934006, -100.93378, -100.93355, -100.93333, -100.93311, -100.9329, -100.932686, -100.93249, -100.93228, -100.93209, -100.93189, -100.9317, -100.93152, -100.93133, -100.931145, -100.930954, -100.93077, -100.93058, -100.9304, -100.93021, -100.93002, -100.92983, -100.92965, -100.92946, -100.929276, -100.92909, -100.92892, -100.928734, -100.928566, -100.92839, -100.92823, -100.92807, -100.92791, -100.927765, -100.92761, -100.927475, -100.92733, -100.9272, -100.92706, -100.926926, -100.926796, -100.92664, -100.92651, -100.92638, -100.92623, -100.92609, -100.92594, -100.9258, -100.925644, -100.92549, -100.92533, -100.92517, -100.92501, -100.92484, -100.92468, -100.924515, -100.92435, -100.92419, -100.92402, -100.92385, -100.92369, -100.92353, -100.92336, -100.9232, -100.92304, -100.92288, -100.92272, -100.92257, -100.92241, -100.92225, -100.9221, -100.921936, -100.92178, -100.92162, -100.92147, -100.92131, -100.92116, -100.921, -100.920845, -100.92069, -100.92053, -100.92038, -100.92023, -100.92007, -100.919914, -100.91976, -100.9196, -100.91945, -100.91929, -100.919136, -100.918976, -100.91882, -100.91866, -100.91859, -100.918434, -100.918274, -100.91812, -100.91797, -100.917816, -100.91767, -100.91753, -100.91738, -100.91724, -100.9171, -100.91696, -100.91683, -100.916695, -100.916565, -100.916435, -100.916306, -100.916176, -100.916046, -100.91592, -100.91579, -100.91566, -100.91553, -100.91539, -100.91525, -100.915115, -100.91498, -100.91483, -100.91469, -100.914536, -100.91439, -100.91424, -100.914085, -100.91393, -100.91377, -100.91362, -100.91346, -100.9133, -100.91314, -100.91298, -100.91282, -100.91266, -100.91249, -100.91232, -100.912155, -100.91198, -100.911804, -100.91163, -100.911446, -100.91126, -100.91106, -100.91087, -100.91068, -100.910484, -100.910286, -100.91009, -100.90988, -100.90968, -100.90948, -100.90927, -100.90906, -100.90885, -100.908646, -100.90843, -100.908226, -100.90801, -100.90781, -100.90759, -100.90739, -100.90717, -100.90696, -100.906746, -100.90653, -100.90632, -100.9061, -100.905876, -100.905655, -100.905426, -100.9052, -100.90497, -100.90473, -100.904495, -100.90426, -100.90402, -100.90378, -100.903534, -100.90329, -100.903046, -100.90281, -100.902565, -100.90232, -100.902084, -100.90184, -100.9016, -100.901375, -100.90114, -100.90091, -100.90068, -100.90045, -100.90022, -100.9, -100.89977, -100.89955, -100.89933, -100.8991, -100.89888, -100.89865, -100.89842, -100.8982, -100.897964, -100.897736, -100.8975, -100.89726, -100.897026, -100.89679, -100.896545, -100.89631, -100.896065, -100.89582, -100.89558, -100.895325, -100.89508, -100.89484, -100.894585, -100.89434, -100.8941, -100.893845, -100.8936, -100.89336, -100.893105, -100.89286, -100.89262, -100.89237, -100.89213, -100.891884, -100.89164, -100.891396, -100.89116, -100.890915, -100.89067, -100.89043, -100.89018, -100.88994, -100.889694, -100.88944, -100.8892, -100.888954, -100.8887, -100.88845, -100.88821, -100.887955, -100.8877, -100.88743, -100.88718, -100.886925, -100.88667, -100.88642, -100.88617, -100.885925, -100.88567, -100.88543, -100.885185, -100.88494, -100.8847, -100.88445, -100.88421, -100.88397, -100.88373, -100.88349, -100.883255, -100.88302, -100.88278, -100.882545, -100.88231, -100.88207, -100.881836, -100.8816, -100.881355, -100.88112, -100.88088, -100.880646, -100.8804, -100.880165, -100.87992, -100.87968, -100.87944, -100.879196, -100.87895, -100.87871, -100.878456, -100.87821, -100.87797, -100.87772, -100.8776, -100.87735, -100.877106, -100.87686, -100.87662, -100.87637, -100.87613, -100.87589, -100.87565, -100.87541, -100.87517, -100.87493, -100.874695, -100.87446, -100.87422, -100.87398, -100.87374, -100.873505, -100.87327, -100.873024, -100.87278, -100.87254, -100.8723, -100.872055, -100.8718, -100.87156, -100.871315, -100.87106, -100.87081, -100.87057, -100.870316, -100.87007, -100.86983, -100.869576, -100.86933, -100.86909, -100.86885, -100.868614, -100.86838, -100.86814, -100.86791, -100.867676, -100.86745, -100.867226, -100.867, -100.866776, -100.866554, -100.86633, -100.86611, -100.86589, -100.86566, -100.86544, -100.86522, -100.86499, -100.86477, -100.86454, -100.86431, -100.86408, -100.86385, -100.863625, -100.863396, -100.86317, -100.86293, -100.8627, -100.86247, -100.86224, -100.86202, -100.86179, -100.86157, -100.86135, -100.86113, -100.860916, -100.86068, -100.860466, -100.86025, -100.86005, -100.85983, -100.85963, -100.85942, -100.859215, -100.85901, -100.8588, -100.8586, -100.8584, -100.85819, -100.85799, -100.85779, -100.85758, -100.857376, -100.85718, -100.85698, -100.85678, -100.85658, -100.85648, -100.856285, -100.856094, -100.8559, -100.85572, -100.85553, -100.85535, -100.85516, -100.85499, -100.854805, -100.85463, -100.854454, -100.85428, -100.854095, -100.85392, -100.85374, -100.85356, -100.85337, -100.85319, -100.853, -100.852806, -100.85261, -100.85241, -100.8522, -100.852, -100.85179, -100.851585, -100.85137, -100.85116, -100.85095, -100.85074, -100.85053, -100.85033, -100.85012, -100.849915, -100.84972, -100.84952, -100.84933, -100.84913, -100.848946, -100.848755, -100.848564, -100.84837, -100.84819, -100.848, -100.84781, -100.84761, -100.84742, -100.84721, -100.847015, -100.84681, -100.846596, -100.84638, -100.84616, -100.84595, -100.84572, -100.8455, -100.84527, -100.84505, -100.84482, -100.8446, -100.844376, -100.844154, -100.84394, -100.84372, -100.84351, -100.8433, -100.843094, -100.84289, -100.84269, -100.84249, -100.84229, -100.842094, -100.841896, -100.8417, -100.84151, -100.84131, -100.84111, -100.84091, -100.84071, -100.840515, -100.84032, -100.8402, -100.840004, -100.839806, -100.83961, -100.83941, -100.83922, -100.83902, -100.83883, -100.83864, -100.83845, -100.83826, -100.83807, -100.83788, -100.8377, -100.83752, -100.83733, -100.83716, -100.836975, -100.83679, -100.83662, -100.83643, -100.83625, -100.836075, -100.83589, -100.83571, -100.835526, -100.83534, -100.83515, -100.83497, -100.83478, -100.834595, -100.834404, -100.83421, -100.83402, -100.83384, -100.83365, -100.83346, -100.83327, -100.833084, -100.83289, -100.83271, -100.83252, -100.83234, -100.83215, -100.83197, -100.83178, -100.8316, -100.83141, -100.83123, -100.83105, -100.83086, -100.83067, -100.83049, -100.8303, -100.83012, -100.829926, -100.82974, -100.82955, -100.82936, -100.82917, -100.82899, -100.8288, -100.828606, -100.82842, -100.82823, -100.82805, -100.82786, -100.827675, -100.82749, -100.82731, -100.82712, -100.82694, -100.82676, -100.82658, -100.82639, -100.82622, -100.826035, -100.82586, -100.825676, -100.8255, -100.825325, -100.82514, -100.82506, -100.824875, -100.8247, -100.824524, -100.82434, -100.824165, -100.82398, -100.82381, -100.82362, -100.82344, -100.82324, -100.82306, -100.822876, -100.82269, -100.82251, -100.82232, -100.822136, -100.82195, -100.82176, -100.82158, -100.821396, -100.821205, -100.821014, -100.82083, -100.82064, -100.82046, -100.82027, -100.82008, -100.81989, -100.81971, -100.81952, -100.819336, -100.81915, -100.81897, -100.81878, -100.818596, -100.81841, -100.81824, -100.818054, -100.81788, -100.817696, -100.81752, -100.817345, -100.81717, -100.817, -100.816826, -100.81666, -100.81649, -100.81632, -100.816154, -100.815994, -100.815834, -100.81567, -100.815506, -100.815346, -100.815186, -100.81503, -100.81487, -100.81471, -100.81455, -100.81439, -100.81431, -100.81415, -100.81398, -100.81381, -100.81365, -100.813484, -100.81331, -100.81314, -100.81297, -100.8128, -100.81262, -100.812454, -100.81228, -100.81211, -100.811935, -100.81177, -100.8116, -100.81143, -100.811264, -100.8111, -100.810936, -100.81077, -100.81061, -100.81044, -100.81028, -100.81012, -100.80996, -100.8098, -100.80964, -100.80948, -100.80932, -100.80916, -100.809006, -100.808846, -100.808685, -100.80853, -100.80838, -100.80822, -100.80807, -100.807915, -100.80777, -100.80762, -100.80755, -100.807396, -100.80725, -100.807106, -100.80696, -100.80682, -100.80668, -100.80653, -100.80639, -100.806244, -100.80608, -100.80594, -100.805786, -100.80564, -100.80549, -100.80534, -100.80519, -100.80504, -100.804886, -100.80473, -100.80458, -100.804436, -100.80428, -100.80413, -100.803986, -100.80384, -100.8037, -100.80356, -100.80342, -100.80328, -100.803154, -100.803024, -100.802895, -100.80277, -100.80265, -100.802536, -100.802414, -100.80231, -100.80219, -100.802086, -100.80198, -100.80187, -100.801765, -100.80167, -100.80156, -100.80146, -100.80136, -100.80126, -100.80116, -100.80106, -100.800964, -100.80087, -100.80077, -100.800674, -100.80058, -100.80048, -100.80039, -100.80029, -100.8002, -100.80011, -100.80002, -100.79992, -100.79983, -100.799736, -100.799644, -100.79955, -100.79946, -100.79937, -100.79928, -100.79918, -100.79909, -100.798996, -100.798904, -100.798805, -100.79871, -100.798615, -100.798515, -100.79842, -100.798325, -100.798225, -100.79813, -100.79803, -100.79792, -100.79782, -100.79772, -100.797615, -100.797516, -100.79741, -100.7973, -100.797195, -100.79709, -100.79698, -100.796875, -100.79676, -100.79665, -100.79654, -100.79643, -100.79632, -100.7962, -100.7961, -100.79598, -100.795876, -100.79582, -100.795715, -100.79561, -100.7955, -100.795395, -100.79529, -100.79519, -100.79508, -100.79498, -100.79488, -100.79477, -100.79467, -100.79457, -100.79447, -100.79437, -100.79427, -100.794174, -100.794075, -100.793976, -100.79388, -100.79378, -100.79368, -100.79358, -100.79348, -100.79338, -100.793274, -100.793175, -100.793076, -100.79298, -100.79288, -100.79278, -100.79267, -100.79257, -100.792465, -100.79236, -100.79226, -100.79215, -100.79204, -100.79193, -100.791824, -100.79171, -100.791595, -100.79148, -100.79137, -100.791245, -100.79112, -100.79101, -100.790886, -100.79076, -100.790634, -100.790504, -100.79038, -100.79025, -100.79012, -100.78999, -100.78986, -100.789734, -100.7896, -100.78947, -100.78933, -100.7892, -100.78906, -100.788925, -100.788795, -100.78866, -100.78852, -100.78838, -100.78825, -100.78812, -100.78798, -100.78784, -100.78771, -100.787575, -100.78744, -100.7873, -100.78716, -100.787025, -100.78689, -100.78675, -100.786606, -100.78647, -100.78632, -100.786255, -100.78611, -100.785965, -100.78581, -100.78567, -100.78552, -100.78537, -100.785225, -100.78507, -100.78492, -100.784775, -100.78462, -100.78447, -100.78432, -100.784164, -100.78401, -100.78385, -100.7837, -100.78354, -100.78337, -100.78321, -100.78304, -100.78287, -100.78269, -100.78252, -100.78233, -100.78215, -100.78196, -100.78177, -100.78158, -100.78138, -100.78118, -100.78098, -100.780785, -100.78058, -100.78038, -100.78018, -100.77998, -100.77978, -100.77958, -100.77939, -100.77917, -100.77898, -100.77878, -100.77859, -100.7784, -100.778206, -100.77802, -100.77783, -100.77765, -100.777466, -100.77728, -100.77709, -100.77691, -100.776726, -100.776535, -100.776344, -100.77615, -100.775955, -100.77576, -100.77555, -100.775345, -100.77514, -100.774925, -100.774704, -100.77448, -100.774254, -100.774025, -100.77379, -100.77355, -100.773315, -100.77307, -100.77283, -100.77258, -100.77234, -100.772095, -100.77186, -100.771614, -100.77137, -100.77113, -100.770905, -100.77067, -100.77044, -100.77021, -100.76999, -100.76977, -100.769554, -100.76933, -100.76912, -100.768906, -100.76869, -100.768486, -100.76827, -100.76806, -100.76784, -100.767624, -100.7674, -100.76718, -100.76696, -100.76673, -100.76651, -100.76627, -100.766045, -100.76581, -100.76557, -100.765335, -100.7651, -100.76486, -100.764626, -100.76439, -100.76415, -100.763916, -100.76368, -100.76344, -100.76321, -100.76298, -100.76274, -100.76251, -100.762276, -100.76205, -100.76182, -100.76159, -100.76137, -100.76114, -100.760925, -100.760704, -100.76049, -100.76028, -100.76007, -100.759865, -100.75967, -100.75947, -100.75928, -100.75908, -100.758896, -100.758705, -100.758514, -100.75833, -100.75815, -100.75796, -100.75777, -100.75758, -100.75739, -100.75718, -100.75698, -100.75678, -100.75658, -100.75637, -100.75616, -100.75595, -100.75573, -100.755516, -100.755295, -100.75507, -100.754845, -100.75462, -100.754395, -100.754166, -100.75394, -100.75371, -100.75349, -100.753265, -100.75304, -100.75282, -100.7526, -100.75239, -100.752174, -100.75197, -100.751755, -100.75155, -100.75135, -100.751144, -100.75094, -100.75074, -100.750534, -100.75033, -100.75012, -100.749916, -100.7497, -100.74948, -100.74926, -100.74904, -100.74881, -100.74857, -100.74834, -100.74809, -100.74785, -100.7476, -100.747345, -100.747086, -100.74683, -100.746574, -100.746315, -100.746056, -100.7458, -100.745544, -100.745285, -100.745026, -100.744774, -100.74452, -100.74428, -100.744026, -100.743774, -100.74353, -100.74328, -100.743034, -100.74278, -100.74253, -100.74228, -100.74203, -100.74177, -100.74151, -100.74125, -100.74098, -100.740715, -100.74045, -100.74032, -100.74004, -100.73977, -100.7395, -100.73923, -100.73895, -100.73868, -100.7384, -100.73814, -100.73786, -100.737724, -100.73746, -100.73718, -100.736916, -100.73665, -100.73638, -100.736115, -100.73585, -100.73558, -100.73532, -100.73502, -100.734764, -100.7345, -100.73424, -100.73397, -100.7337, -100.73344, -100.73317, -100.7329, -100.73263, -100.73236, -100.73208, -100.731804, -100.73152, -100.73124, -100.73095, -100.73066, -100.73037, -100.73007, -100.729774, -100.72963, -100.729324, -100.72902, -100.728714, -100.72841, -100.7281, -100.7278, -100.72749, -100.72719, -100.72689, -100.726585, -100.72643, -100.726135, -100.72584, -100.72554, -100.72524, -100.72495, -100.724655, -100.724365, -100.72407, -100.72378, -100.72348, -100.723335, -100.72304, -100.72274, -100.72244, -100.722145, -100.72185, -100.72155, -100.72125, -100.720955, -100.72066, -100.72036, -100.72006, -100.71977, -100.71948, -100.71919, -100.71891, -100.71863, -100.718346, -100.71807, -100.7178, -100.71752, -100.717255, -100.71698, -100.71671, -100.716446, -100.71618, -100.715904, -100.71564, -100.71536, -100.71509, -100.71481, -100.71453, -100.71426, -100.713974, -100.713684, -100.7134, -100.71311, -100.71282, -100.71253, -100.71224, -100.71196, -100.71167, -100.711525, -100.711235, -100.710945, -100.710655, -100.71037, -100.71008, -100.70979, -100.70951, -100.70922, -100.70893, -100.708786, -100.708496, -100.708206, -100.70792, -100.70762, -100.70733, -100.70703, -100.706726, -100.70643, -100.70612, -100.705826, -100.70567, -100.70537, -100.70506, -100.70476, -100.704445, -100.70414, -100.70383, -100.703514, -100.7032, -100.70305, -100.70273, -100.70254, -100.70222, -100.7019, -100.70158, -100.701256, -100.700935, -100.700615, -100.700294, -100.699974, -100.69965, -100.69934, -100.69903, -100.698715, -100.69841, -100.698105, -100.69781, -100.69751, -100.69722, -100.69694, -100.69665, -100.69637, -100.6961, -100.69582, -100.69555, -100.69528, -100.695015, -100.69475, -100.69448, -100.69422, -100.69396, -100.6937, -100.693565, -100.693306, -100.69305, -100.69279, -100.69253, -100.69227, -100.69201, -100.69175, -100.69148, -100.69122, -100.690956, -100.69068, -100.690414, -100.69014, -100.689865, -100.68959, -100.68931, -100.689026, -100.68874, -100.68846, -100.68817, -100.68789, -100.6876, -100.68732, -100.68703, -100.686745, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -100.63909, -100.63877, -100.63845, -100.63813, -100.63781, -100.63749, -100.63716, -100.63684, -100.63651, -100.63619, -100.635864, -100.635544, -100.635216, -100.634895, -100.63457, -100.63425, -100.63392, -100.6336, -100.63328, -100.63295, -100.63263, -100.63231, -100.63198, -100.63166, -100.63134, -100.63102, -100.63069, -100.63037, -100.63004, -100.62972, -100.629395, -100.62907, -100.62874, -100.62841, -100.628075, -100.62775, -100.62741, -100.627075, -100.62674, -100.6264, -100.62607, -100.625725, -100.62556, -100.62522, -100.624886, -100.62455, -100.62421, -100.62387, -100.623535, -100.6232, -100.62286, -100.62253, -100.622185, -100.62185, -100.62151, -100.62118, -100.62084, -100.62051, -100.62016, -100.61983, -100.619484, -100.61915, -100.618805, -100.61863, -100.618286, -100.61794, -100.6176, -100.617256, -100.616905, -100.61656, -100.61622, -100.61587, -100.615524, -100.61517, -100.61483, -100.61448, -100.61413, -100.613785, -100.613434, -100.61308, -100.61273, -100.61238, -100.61203, -100.61168, -100.61133, -100.61098, -100.61062, -100.61027, -100.60991, -100.60956, -100.6092, -100.60885, -100.60849, -100.6081, -100.60774, -100.60738, -100.60703, -100.606674, -100.60632, -100.605965, -100.60561, -100.605255, -100.604904, -100.60455, -100.6042, -100.60385, -100.6035, -100.60315, -100.602806, -100.602455, -100.60211, -100.60176, -100.60142, -100.601074, -100.60073, -100.600555, -100.60021, -100.59987, -100.59952, -100.59917, -100.598816, -100.598465, -100.598114, -100.597755, -100.5974, -100.59704, -100.59668, -100.59632, -100.595955, -100.5956, -100.59523, -100.594864, -100.594505, -100.59414, -100.59377, -100.593414, -100.59305, -100.59268, -100.59232, -100.59196, -100.5916, -100.59124, -100.59088, -100.59052, -100.590164, -100.58981, -100.58946, -100.58929, -100.588936, -100.588585, -100.58824, -100.5879, -100.587555, -100.58721, -100.58687, -100.586525, -100.58636, -100.58601, -100.58567, -100.58532, -100.58498, -100.584625, -100.584274, -100.583916, -100.58356, -100.5832, -100.58284, -100.58266, -100.58229, -100.581924, -100.58155, -100.581184, -100.58082, -100.580444, -100.58008, -100.57971, -100.579346, -100.57899, -100.578804, -100.57845, -100.578094, -100.57775, -100.5774, -100.57706, -100.57671, -100.57638, -100.57604, -100.575676, -100.57534, -100.575005, -100.57467, -100.57433, -100.574, -100.573654, -100.57332, -100.572975, -100.57263, -100.57229, -100.571945, -100.57177, -100.57143, -100.571075, -100.57073, -100.57038, -100.57004, -100.56969, -100.56934, -100.56899, -100.56865, -100.568306, -100.56814, -100.567795, -100.56745, -100.567116, -100.56678, -100.566444, -100.56611, -100.56577, -100.565445, -100.56511, -100.56478, -100.56461, -100.564285, -100.56396, -100.56363, -100.5633, -100.56297, -100.562645, -100.56231, -100.56197, -100.561646, -100.56148, -100.56114, -100.56081, -100.56046, -100.56013, -100.559784, -100.55944, -100.559105, -100.55876, -100.55842, -100.558075, -100.55773, -100.55738, -100.55704, -100.556694, -100.55635, -100.55601, -100.55567, -100.55533, -100.554985, -100.55464, -100.554474, -100.55413, -100.55379, -100.553444, -100.5531, -100.55275, -100.55241, -100.552055, -100.551704, -100.55135, -100.551, -100.550644, -100.550285, -100.54992, -100.54956, -100.549194, -100.54882, -100.548454, -100.54809, -100.547714, -100.54734, -100.546974, -100.5466, -100.546234, -100.54587, -100.54551, -100.54514, -100.544785, -100.54443, -100.54408, -100.54373, -100.543564, -100.54322, -100.54288, -100.54254, -100.542206, -100.54187, -100.54153, -100.54119, -100.540855, -100.54051, -100.540344, -100.53999, -100.53965, -100.5393, -100.53895, -100.5386, -100.53824, -100.53788, -100.53752, -100.537155, -100.53676, -100.53639, -100.53603, -100.53567, -100.5353, -100.534935, -100.53457, -100.5342, -100.53384, -100.53347, -100.533104, -100.53292, -100.532555, -100.53218, -100.53181, -100.53143, -100.53106, -100.530685, -100.53031, -100.52993, -100.52956, -100.529175, -100.528984, -100.5286, -100.52822, -100.52784, -100.52746, -100.52708, -100.52669, -100.526306, -100.52592, -100.525536, -100.52515, -100.52495, -100.52456, -100.52417, -100.52377, -100.523384, -100.52298, -100.52258, -100.52218, -100.52177, -100.52136, -100.52095, -100.52074, -100.520325, -100.5199, -100.51948, -100.51905, -100.518616, -100.51819, -100.51775, -100.51733, -100.51689, -100.51646, -100.51624, -100.515816, -100.51538, -100.51495, -100.51453, -100.5141, -100.51368, -100.51325, -100.51283, -100.51241, -100.51199, -100.51157, -100.51116, -100.51074, -100.51032, -100.50991, -100.50949, -100.50907, -100.50865, -100.508224, -100.507805, -100.507385, -100.50696, -100.50653, -100.5061, -100.50568, -100.50524, -100.504814, -100.50438, -100.503944, -100.50351, -100.503296, -100.50286, -100.50242, -100.50198, -100.50155, -100.50111, -100.50067, -100.50023, -100.499794, -100.49931, -100.49887, -100.49843, -100.49799, -100.49755, -100.497116, -100.49667, -100.49624, -100.4958, -100.49536, -100.49493, -100.494705, -100.49427, -100.49383, -100.49339, -100.49295, -100.492516, -100.49207, -100.49163, -100.49119, -100.490746, -100.4903, -100.48985, -100.48941, -100.48896, -100.48851, -100.48806, -100.48761, -100.48715, -100.4867, -100.48625, -100.485794, -100.48557, -100.485115, -100.484665, -100.48421, -100.48376, -100.4833, -100.48285, -100.48239, -100.48194, -100.48148, -100.481255, -100.4808, -100.48034, -100.47988, -100.479416, -100.47896, -100.47849, -100.478035, -100.47757, -100.477104, -100.47664, -100.47617, -100.47594, -100.47547, -100.475006, -100.47453, -100.47407, -100.4736, -100.47314, -100.472664, -100.4722, -100.47173, -100.47127, -100.470795, -100.47033, -100.46986, -100.46939, -100.46892, -100.468445, -100.46797, -100.4675, -100.467026, -100.46678, -100.4663, -100.46582, -100.46534, -100.46486, -100.46437, -100.46388, -100.463394, -100.46291, -100.462425, -100.46194, -100.46145, -100.46121, -100.460724, -100.46024, -100.45976, -100.45928, -100.4588, -100.45832, -100.45785, -100.457375, -100.4569, -100.45643, -100.455956, -100.45548, -100.45501, -100.45454, -100.45406, -100.45359, -100.45312, -100.45264, -100.45216, -100.45187, -100.4514, -100.45092, -100.45044, -100.44996, -100.44948, -100.449, -100.44852, -100.44804, -100.44755, -100.44731, -100.44682, -100.44634, -100.44586, -100.44538, -100.4449, -100.44442, -100.44394, -100.44346, -100.44298, -100.442505, -100.442024, -100.44154, -100.44106, -100.44058, -100.4401, -100.43962, -100.43914, -100.43865, -100.43817, -100.43769, -100.43745, -100.436966, -100.436485, -100.436, -100.43552, -100.435036, -100.434555, -100.434074, -100.43359, -100.43311, -100.43263, -100.43216, -100.43169, -100.43121, -100.43074, -100.43027, -100.42979, -100.429306, -100.428825, -100.428345, -100.427864, -100.42739, -100.42693, -100.42652, -100.42617, -100.42589, -100.42567, -100.425514, -100.42543, -100.4254, -100.42539, -100.4254, -100.425415, -100.425415, -100.42543, -100.42544, -100.425446, -999.0}
alt =
  {955.1, -999.0, -999.0, -999.0, -999.0, -999.0, 956.80334, 960.42993, 964.12164, 967.88635, 971.7343, 975.67664, 979.72455, 983.8871, 988.1648, 992.5561, 997.0593, 1001.67145, 1006.38306, 1011.1833, 1016.0612, 1021.006, 1026.0082, 1031.0587, 1036.1484, 1041.2678, 1046.4064, 1051.5533, 1056.6979, 1061.8295, 1066.9385, 1072.0153, 1077.0505, 1082.035, 1086.9594, 1091.8143, 1096.5912, 1101.2808, 1105.8761, 1110.3707, 1114.7579, 1119.0323, 1123.194, 1127.2441, 1131.1844, 1135.0168, 1138.7451, 1142.3734, 1145.906, 1149.3472, 1152.6998, 1155.967, 1159.1516, 1162.2572, 1165.2922, 1168.2664, 1171.1891, 1174.0696, 1176.9144, 1179.729, 1182.7968, 1185.5641, 1188.3069, 1191.0192, 1193.6951, 1196.3298, 1198.9224, 1201.4727, 1203.9807, 1206.4462, 1208.8691, 1211.2494, 1213.5867, 1215.8785, 1218.1141, 1220.2802, 1222.3634, 1224.3507, 1226.2288, 1227.9846, 1229.6051, 1231.0782, 1232.3966, 1233.5535, 1234.5427, 1235.3606, 1236.015, 1236.5167, 1236.8766, 1237.1077, 1237.2312, 1237.271, -999.0, -999.0, -999.0, -999.0, -999.0, 1237.4781, 1237.8883, 1238.5198, 1239.4148, 1240.612, 1242.1316, 1243.9886, 1246.1984, 1248.7725, 1251.7057, 1254.9883, 1258.6105, 1262.5602, 1266.8156, 1271.3514, 1276.1433, 1281.1658, 1286.3926, 1291.797, 1297.3523, 1303.0311, 1308.8031, 1314.6371, 1320.5021, 1326.3678, 1332.2096, 1338.0048, 1343.73, 1349.3641, 1354.8938, 1360.3086, 1365.5977, 1370.7506, 1375.7579, 1380.6106, 1385.2993, 1389.8164, 1394.1606, 1398.3331, 1402.3348, 1406.1677, 1409.8376, 1413.3522, 1416.7186, 1419.945, 1423.0419, 1426.0209, 1428.8938, 1431.6732, 1434.3787, 1437.0315, 1439.6534, 1442.2651, 1444.8844, 1447.5275, 1450.2109, 1452.95, 1455.7522, 1458.6229, 1461.5676, 1464.59, 1467.6853, 1471.1658, 1474.3903, 1477.6635, 1480.9716, 1484.2997, 1487.633, 1490.9583, 1494.2699, 1497.5643, 1500.8379, 1504.0885, 1507.3203, 1510.539, 1513.7502, 1516.9603, 1520.177, 1523.4084, 1526.6627, 1529.9478, 1533.2697, 1536.6339, 1540.0461, 1543.5118, 1547.0374, 1550.6287, 1554.292, 1558.0338, 1561.8623, 1565.786, 1569.8134, 1573.9519, 1578.2046, 1582.5731, 1587.059, 1591.6611, 1596.3663, 1601.1575, 1606.0176, 1610.9286, 1615.8687, 1620.8147, 1625.7434, 1630.6328, 1635.4672, 1640.2323, 1644.9143, 1649.4998, 1653.979, 1658.3436, 1662.5851, 1666.6959, 1670.6725, 1674.5128, 1678.215, 1681.7782, 1685.2104, 1688.5221, 1691.7236, 1694.8264, 1697.8469, 1700.8035, 1703.7142, 1706.5966, 1709.4637, 1712.3278, 1715.2004, 1718.0927, 1721.0098, 1723.9552, 1726.9326, 1729.9448, 1732.9922, 1736.0739, 1739.1891, 1742.3362, 1745.5099, 1748.7029, 1751.9084, 1755.119, 1758.3262, 1761.5206, 1764.6931, 1767.8342, 1770.9331, 1773.9784, 1776.9585, 1779.8632, 1782.6874, 1785.4282, 1788.0828, 1790.649, 1793.1306, 1795.5331, 1797.8618, 1800.1232, 1802.3251, 1804.477, 1806.5884, 1808.6683, 1810.7262, 1812.7712, 1814.8131, 1816.8604, 1818.9188, 1821.2014, 1823.298, 1825.4183, 1827.5588, 1829.7144, 1831.8794, 1834.0476, 1836.2075, 1838.3463, 1840.451, 1842.5093, 1844.5104, 1846.445, 1848.3031, 1850.0757, 1851.7559, 1853.3374, 1854.8145, 1856.1807, 1857.4298, 1858.5554, 1859.551, 1860.4105, 1861.13, 1861.706, 1862.135, 1862.4147, 1862.5469, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 1863.2009, 1865.7286, 1868.3383, 1871.04, 1873.8473, 1876.7739, 1879.8345, 1883.3721, 1886.7552, 1890.3077, 1894.0393, 1897.9589, 1902.0697, 1906.3735, 1910.8721, 1915.5659, 1920.4495, 1925.5149, 1930.7545, 1936.1598, 1941.7191, 1947.4193, 1953.2473, 1959.1895, 1965.2278, 1971.3436, 1977.5176, 1983.7307, 1989.963, 1996.1941, 2002.4038, 2008.572, 2014.6814, 2020.7152, 2026.6565, 2032.4893, 2038.2017, 2043.7834, 2049.2244, 2054.5154, 2059.6567, 2064.6511, 2069.5022, 2074.2134, 2078.7893, 2083.2358, 2087.5583, 2091.763, 2095.858, 2099.8528, 2103.7573, 2107.5808, 2111.3337, 2115.026, 2118.6677, 2122.2695, 2125.8398, 2129.3867, 2132.9177, 2136.4414, 2139.9631, 2143.4888, 2147.0237, 2150.5725, 2154.1384, 2157.723, 2161.328, 2164.9543, 2168.6006, 2172.2634, 2175.9392, 2179.6255, 2183.323, 2187.0344, 2190.762, 2194.5085, 2198.2817, 2202.0908, 2205.945, 2209.8538, 2213.8274, 2217.8767, 2222.0122, 2226.245, 2230.587, 2235.0493, 2239.6448, 2244.3843, 2249.2764, 2254.3274, 2259.5435, 2264.931, 2270.4902, 2276.2207, 2282.121, 2288.1897, 2294.4192, 2300.8003, 2307.3237, 2314.6523, 2321.4448, 2328.353, 2335.3687, 2342.484, 2349.6887, 2356.973, 2364.3262, 2371.738, 2379.1948, 2386.6829, 2394.188, 2401.696, 2409.194, 2416.6692, 2424.1086, 2431.5002, 2438.8384, 2446.1187, 2453.338, 2460.493, 2467.585, 2474.6172, 2481.5928, 2488.5156, 2495.3938, 2502.237, 2509.0557, 2515.8586, 2522.6506, 2529.434, 2536.2117, 2542.9858, 2549.7554, 2556.5183, 2563.272, 2570.0146, 2576.747, 2583.4707, 2590.1877, 2596.8997, 2603.608, 2610.3132, 2617.017, 2623.7207, 2630.4246, 2637.1294, 2643.8362, 2650.5454, 2657.256, 2663.9668, 2670.676, 2677.3823, 2684.082, 2690.771, 2697.445, 2704.0999, 2710.733, 2717.3416, 2723.9236, 2730.477, 2737.0051, 2743.5122, 2750.0032, 2756.4836, 2762.9617, 2769.4465, 2775.948, 2782.476, 2789.041, 2795.6548, 2802.3286, 2809.0732, 2815.894, 2822.7935, 2829.7742, 2836.8386, 2843.9836, 2851.204, 2858.495, 2865.8503, 2873.2563, 2880.6953, 2888.1504, 2895.6038, 2903.038, 2910.436, 2917.7798, 2925.0525, 2932.2402, 2939.3315, 2946.3147, 2953.1785, 2959.9202, 2966.541, 2973.0427, 2979.4277, 2985.7087, 2991.9038, 2998.0308, 3004.1077, 3010.151, 3016.1763, 3022.1992, 3028.2349, 3034.293, 3040.3801, 3046.5024, 3052.6665, 3058.871, 3065.1123, 3071.3855, 3078.3167, 3084.6296, 3090.934, 3097.2107, 3103.4402, 3109.6028, 3115.679, 3121.649, 3127.4937, 3133.202, 3138.7642, 3144.172, -999.0, -999.0, -999.0, 3164.2385, 3168.901, 3173.4385, 3177.8596, 3182.1729, 3186.387, 3190.5076, 3194.5398, 3198.4888, 3202.359, 3206.1533, 3209.8733, 3213.5208, 3217.0972, 3220.602, 3224.0344, 3227.393, 3230.677, 3233.885, 3237.017, 3240.0728, 3243.0515, 3245.9563, 3248.7908, 3251.5586, 3254.2637, 3256.915, 3259.5225, 3262.0964, 3264.6472, 3267.1865, 3269.7258, 3272.2769, 3274.8518, 3277.463, 3280.1223, 3282.8425, 3285.6353, 3288.5073, 3291.4626, 3294.5051, 3297.638, 3300.856, 3304.1506, 3307.5125, 3310.933, 3314.4084, 3317.9363, 3321.5151, 3325.1436, 3328.8252, 3332.5664, 3336.3735, 3340.253, 3344.2078, 3348.2397, 3352.351, 3356.5422, 3360.8054, 3365.127, 3369.4934, 3373.8914, 3378.3062, 3382.7224, 3387.125, 3391.4993, 3395.8354, 3400.1272, 3404.3687, 3408.5535, 3412.6787, 3416.7441, 3420.7483, 3424.6907, 3428.5713, 3432.3904, 3436.1484, 3440.2117, 3443.8418, 3447.4111, 3450.9197, 3454.3682, 3457.7642, 3461.1177, 3464.4392, 3467.7393, 3471.0317, 3474.3318, 3477.6553, 3481.0164, 3484.425, 3487.8892, 3491.4163, 3495.013, 3498.6807, 3502.4182, 3506.224, 3510.0964, 3514.0298, 3518.0168, 3522.0505, 3526.1235, 3530.2278, 3534.356, 3538.4995, 3542.6516, 3546.8096, 3550.9739, 3555.145, 3559.323, 3563.5105, 3567.7107, 3571.9268, 3576.1616, 3580.417, 3584.6929, 3588.99, 3593.3093, 3597.6543, 3602.0315, 3606.4463, 3610.9045, 3615.414, 3619.9827, 3624.6182, 3629.328, 3634.1086, 3638.9521, 3643.8499, 3648.793, 3653.7715, 3658.7737, 3663.7878, 3668.8037, 3673.8203, 3678.8416, 3683.8713, 3688.9143, 3693.977, 3699.0676, 3704.1938, 3709.3635, 3714.5806, 3719.8477, 3725.1665, 3730.539, 3735.963, 3741.433, 3746.945, 3752.4934, 3758.0688, 3763.6606, 3769.2576, 3774.8484, 3780.4238, 3785.976, 3791.4973, 3796.9792, 3802.4158, 3807.8025, 3813.1343, 3818.4058, 3823.6125, 3828.7493, 3833.8108, 3838.7927, 3843.6934, 3848.5137, 3853.2546, 3857.917, 3862.504, 3867.019, 3871.4666, 3875.8503, 3880.1716, 3884.4304, 3888.627, 3892.7607, 3896.8303, 3901.2292, 3905.1553, 3909.0085, 3912.784, 3916.475, 3920.0757, 3923.579, 3926.9766, 3930.2573, 3933.412, 3936.4307, 3939.3086, 3942.0437, 3944.6335, 3947.0764, 3949.3762, 3951.5396, 3953.5725, 3955.4827, 3957.2793, 3958.9739, 3960.5781, 3962.1035, 3963.5615, 3964.964, 3966.323, 3967.6501, 3968.9575, 3970.258, 3971.5635, 3972.886, 3974.234, 3975.6133, 3977.0298, 3978.4895, 3979.994, 3981.5435, 3983.1377, 3984.7764, 3986.457, 3988.176, 3989.9294, 3991.7134, 3993.5222, 3995.3489, 3997.1868, 3999.0288, 4000.87, 4002.706, 4004.5327, 4006.346, 4008.1453, 4009.0403, 4010.822, 4012.5945, 4014.36, 4016.1245, 4017.893, 4019.6714, 4021.465, 4023.2815, 4025.1274, 4027.0103, 4028.9363, 4030.91, 4032.9355, 4035.0173, 4037.1577, 4039.3547, 4041.6052, 4043.9065, 4046.256, 4048.6523, 4051.0928, 4053.5762, 4056.0999, 4058.6611, 4061.2568, 4063.8833, 4066.539, 4069.2256, 4071.9456, 4074.701, 4077.496, 4080.3394, 4083.2402, 4086.2083, 4089.2532, 4092.387, 4095.6213, 4098.9688, 4102.44, 4106.045, 4109.7925, 4113.6924, 4117.7515, 4121.9697, 4126.347, 4130.8823, 4135.5713, 4140.4, 4145.351, 4150.9194, 4156.074, 4161.2983, 4166.573, 4171.879, 4177.198, 4182.513, 4187.8057, 4193.059, 4198.258, 4203.3896, 4208.444, 4213.4097, 4218.278, 4223.0444, 4227.7065, 4232.261, 4236.7065, 4241.047, 4245.2856, 4249.4272, 4253.477, 4257.4434, 4261.334, 4265.157, 4268.922, 4272.637, 4276.314, 4279.961, 4283.588, 4287.201, 4290.806, 4294.4097, 4298.018, 4301.638, 4305.2764, 4308.94, 4312.6333, 4316.3555, 4320.105, 4323.881, 4327.6797, 4331.498, 4335.332, 4339.177, 4343.0283, 4346.8833, 4350.7373, 4354.587, 4358.43, 4362.267, 4366.099, 4369.9277, 4373.753, 4377.5693, 4381.373, 4385.159, 4388.922, 4392.6543, 4396.349, 4399.9985, 4403.5967, 4407.1387, 4410.62, 4414.037, 4417.386, 4420.665, 4423.8716, 4427.004, 4430.063, 4433.055, 4435.9883, 4438.8696, 4441.7085, 4444.517, 4447.309, 4450.0967, 4452.893, 4455.7075, 4458.55, 4461.429, 4464.3535, 4467.3296, 4470.3623, 4473.458, 4476.6206, 4479.852, 4483.1553, 4486.5312, 4489.9814, 4493.506, 4497.1035, 4500.7734, 4504.5146, 4508.3223, 4512.1904, 4516.114, 4520.087, 4524.1016, 4528.151, 4532.226, 4536.322, 4540.8496, 4544.9863, 4549.1426, 4553.3174, 4557.5073, 4561.708, 4565.915, 4570.1255, 4574.3335, 4578.5347, 4582.724, 4586.8994, 4591.064, 4595.22, 4599.373, 4603.524, 4607.6753, 4611.8267, 4615.9795, 4620.134, 4624.289, 4628.444, 4632.5977, 4636.749, 4640.8975, 4645.041, 4649.1787, 4653.31, 4657.4355, 4661.5576, 4665.6772, 4669.797, 4673.9214, 4678.0547, 4682.202, 4686.367, 4690.553, 4694.7617, 4698.9956, 4703.2554, 4707.538, 4709.6875, 4714.0, 4718.328, 4722.671, 4727.029, 4731.4023, 4735.7915, 4740.195, 4744.6113, 4749.0386, 4753.474, 4757.915, 4762.356, 4766.7925, 4771.2197, 4775.6353, 4780.038, 4784.4272, 4788.8022, 4793.161, 4797.504, 4801.8286, 4806.135, 4810.4214, 4814.6865, 4818.9297, 4823.149, 4827.3457, 4831.523, 4835.6836, 4839.83, 4843.9653, 4848.0913, 4852.21, 4856.323, 4860.4336, 4864.544, 4868.6567, 4872.774, 4876.8994, 4881.0356, 4885.187, 4889.3564, 4893.545, 4897.75, 4901.9717, 4906.2075, 4910.455, 4914.71, 4918.969, 4923.2285, 4927.4844, 4931.735, 4935.976, 4940.2065, 4944.4253, 4948.6353, 4952.838, 4957.0356, 4961.2314, 4965.428, 4969.629, 4973.837, 4978.0576, 4982.2964, 4986.5605, 4990.8564, 4995.19, 4999.569, 5003.9985, 5008.487, 5013.0376, 5018.1196, 5022.812, 5027.576, 5032.4146, 5037.3276, 5042.317, 5047.384, 5052.525, 5057.7373, 5063.016, 5068.3564, 5073.756, 5079.211, 5084.7188, 5090.277, 5095.8833, 5101.5386, 5107.2437, 5112.9976, 5118.7993, 5124.6475, 5127.588, 5133.5005, 5139.4526, 5145.4375, 5151.4478, 5157.4766, 5163.515, 5169.5557, 5175.5874, 5181.601, 5187.588, 5193.5425, 5199.4595, 5205.333, 5211.1587, 5216.9316, 5222.647, 5228.3003, 5233.888, 5239.409, 5244.862, 5250.2456, 5255.561, 5260.813, 5266.006, 5271.146, 5276.2383, 5281.289, 5286.3057, 5291.294, 5296.26, 5301.2026, 5306.122, 5311.018, 5315.8887, 5320.73, 5325.5376, 5330.3066, 5335.033, 5339.7134, 5344.344, 5348.9224, 5353.4453, 5357.9155, 5362.3354, 5366.7075, 5371.0356, 5375.3306, 5379.603, 5383.8647, 5388.1255, 5392.3916, 5396.668, 5400.959, 5405.27, 5409.603, 5413.9585, 5418.3384, 5422.743, 5427.171, 5431.618, 5436.082, 5440.559, 5445.0454, 5449.5366, 5454.028, 5458.5156, 5463.0015, 5467.4863, 5471.973, 5476.4634, 5480.9624, 5485.476, 5490.01, 5494.5684, 5499.1587, 5503.786, 5508.457, 5513.176, 5517.947, 5522.772, 5527.6553, 5530.614, 5535.592, 5540.6255, 5545.712, 5550.848, 5556.0273, 5561.241, 5566.48, 5571.7354, 5576.998, 5582.2607, 5587.5166, 5592.7573, 5597.977, 5603.171, 5608.3345, 5613.463, 5618.552, 5623.598, 5628.599, 5633.5513, 5638.453, 5643.3037, 5648.103, 5652.8506, 5657.5483, 5662.199, 5666.8066, 5671.374, 5675.9043, 5680.401, 5684.867, 5689.306, 5693.7217, 5698.118, 5702.5, 5706.8726, 5711.239, 5715.6025, 5719.968, 5724.3374, 5728.712, 5733.0894, 5737.467, 5741.842, 5746.2104, 5750.5684, 5754.9106, 5759.2324, 5763.5303, 5767.8027, 5772.047, 5776.2617, 5780.4487, 5784.614, 5788.763, 5792.903, 5797.036, 5801.1675, 5805.2993, 5809.4346, 5813.575, 5817.722, 5821.877, 5826.0396, 5830.21, 5834.387, 5838.569, 5842.7544, 5846.94, 5851.1216, 5855.2944, 5859.4536, 5863.597, 5867.7236, 5871.832, 5875.9214, 5879.992, 5884.045, 5888.0815, 5892.1025, 5896.112, 5898.114, 5902.116, 5906.121, 5910.1343, 5914.16, 5918.202, 5922.2637, 5926.349, 5930.4614, 5934.604, 5939.1987, 5943.414, 5947.67, 5951.9697, 5956.3174, 5960.716, 5965.1694, 5969.68, 5974.2515, 5978.8857, 5983.5815, 5988.3394, 5993.157, 5998.0337, 6002.965, 6007.9473, 6012.976, 6018.047, 6023.156, 6028.2983, 6033.4697, 6038.6655, 6043.877, 6049.0957, 6054.314, 6059.522, 6064.7104, 6069.8677, 6074.9834, 6080.05, 6085.065, 6090.0303, 6094.947, 6099.816, 6104.64, 6109.423, 6114.168, 6118.879, 6123.56, 6128.217, 6132.853, 6137.474, 6142.085, 6146.689, 6151.2915, 6155.896, 6160.5093, 6165.1357, 6169.7812, 6174.452, 6179.1543, 6181.519, 6186.2812, 6191.0913, 6195.9565, 6200.883, 6205.8765, 6210.944, 6216.0854, 6221.297, 6226.5728, 6231.9087, 6237.3003, 6242.746, 6248.242, 6253.787, 6259.3784, 6265.0166, 6270.7, 6276.429, 6282.204, 6288.027, 6293.8994, 6299.823, 6305.802, 6311.8374, 6317.935, 6324.0977, 6330.326, 6336.619, 6342.9736, 6349.3877, 6355.8584, 6362.3804, 6368.9487, 6375.558, 6382.204, 6388.8813, 6395.585, 6402.31, 6409.052, 6415.804, 6422.563, 6425.9424, 6432.7, 6439.4517, 6446.193, 6452.921, 6459.6313, 6466.3237, 6472.9976, 6479.6514, 6486.2856, 6493.559, 6500.1484, 6506.715, 6513.2583, 6519.7793, 6526.2783, 6532.757, 6539.216, 6545.6577, 6552.085, 6558.5, 6564.9062, 6571.3105, 6577.7197, 6584.1416, 6590.582, 6597.045, 6603.533, 6610.0493, 6616.596, 6623.1743, 6629.7827, 6636.421, 6643.089, 6649.7837, 6656.503, 6663.2437, 6670.003, 6676.779, 6683.569, 6690.371, 6697.183, 6704.0015, 6710.821, 6717.638, 6724.4497, 6731.2515, 6738.0415, 6744.817, 6751.575, 6758.312, 6765.0234, 6771.706, 6778.3564, 6784.9736, 6791.5576, 6798.109, 6804.627, 6811.113, 6817.5674, 6823.992, 6830.3877, 6836.756, 6843.0977, 6849.416, 6855.712, 6861.988, 6868.247, 6874.4927, 6880.726, 6886.9478, 6893.157, 6899.353, 6905.535, 6911.7026, 6917.8545, 6923.9897, 6930.1074, 6936.2085, 6942.2935, 6948.362, 6954.414, 6960.442, 6966.4375, 6972.3906, 6978.293, 6984.141, 6989.9307, 6995.658, 7001.3213, 7006.917, 7012.4443, 7017.902, 7023.288, 7028.6025, 7033.847, 7039.0215, 7044.1265, 7049.164, 7054.136, 7059.0444, 7063.89, 7066.2905, 7071.046, 7075.741, 7080.3784, 7084.959, 7089.4883, 7093.9697, 7098.408, 7102.808, 7107.172, 7111.9346, 7116.2344, 7120.5093, 7124.765, 7129.0073, 7133.241, 7137.471, 7141.703, 7145.941, 7150.19, 7154.454, 7158.737, 7163.0405, 7167.368, 7171.7227, 7176.107, 7180.523, 7184.9727, 7189.4546, 7193.962, 7198.4873, 7203.0244, 7207.566, 7212.1055, 7216.6357, 7221.151, 7225.645, 7230.1133, 7234.552, 7238.9565, 7243.3228, 7247.645, 7251.9194, 7256.141, 7260.309, 7264.427, 7268.4985, 7272.5273, 7276.5176, 7280.472, 7284.3955, 7288.29, 7292.158, 7295.9995, 7299.8135, 7303.5996, 7307.359, 7311.0947, 7314.8086, 7318.5044, 7322.184, 7325.8506, 7329.505, 7333.1504, 7336.789, 7340.4233, 7344.056, 7347.6895, 7351.3267, 7354.971, 7358.6274, 7362.298, 7365.9893, 7369.7085, 7373.4644, 7377.264, 7381.116, 7385.0283, 7389.01, 7393.068, 7397.2114, 7401.4507, 7403.6094, 7408.01, 7412.53, 7417.1743, 7421.949, 7426.859, 7431.9077, 7437.0967, 7442.425, 7447.892, 7453.497, 7459.239, 7465.1147, 7471.1226, 7477.2607, 7483.523, 7489.904, 7496.396, 7502.9937, 7509.684, 7516.4546, 7523.291, 7530.179, 7537.103, 7544.044, 7550.984, 7557.905, 7564.782, 7571.591, 7578.3057, 7584.9014, 7591.363, 7597.676, 7603.8267, 7609.8047, 7615.6113, 7621.2534, 7626.7383, 7632.0737, 7637.2705, 7642.3423, 7647.793, 7652.6445, 7657.407, 7662.09, 7666.701, 7671.2495, 7675.7427, 7680.1904, 7684.6, 7688.9805, 7693.341, 7697.6895, 7702.035, 7706.3867, 7710.751, 7715.1333, 7719.541, 7723.979, 7728.4478, 7732.947, 7737.475, 7742.0327, 7746.6177, 7751.2305, 7755.869, 7760.5337, 7765.2227, 7769.9346, 7774.6675, 7779.4204, 7784.1943, 7788.99, 7793.8096, 7798.6533, 7803.519, 7808.4033, 7813.3037, 7818.217, 7823.144, 7828.0884, 7833.0513, 7838.035, 7843.0425, 7848.0737, 7853.131, 7858.215, 7863.3257, 7868.463, 7873.625, 7878.8125, 7884.023, 7889.255, 7894.5073, 7899.7773, 7905.0615, 7910.356, 7915.656, 7920.957, 7926.2593, 7931.5625, 7936.867, 7942.1733, 7947.483, 7952.799, 7958.1235, 7963.4585, 7968.8047, 7974.1626, 7979.532, 7984.913, 7990.306, 7995.7114, 8001.129, 8006.56, 8012.0093, 8017.4844, 8022.991, 8028.537, 8034.1304, 8039.7803, 8045.4956, 8051.2847, 8057.1514, 8063.098, 8069.127, 8075.24, 8081.437, 8087.718, 8094.08, 8100.524, 8107.043, 8113.631, 8120.2812, 8126.9863, 8133.7363, 8140.521, 8147.3296, 8154.1514, 8160.977, 8167.7964, 8174.6006, 8181.381, 8188.8013, 8195.505, 8202.16, 8208.761, 8215.298, 8221.764, 8228.151, 8234.453, 8240.658, 8246.759, 8252.744, 8258.605, 8264.333, 8269.915, 8275.343, 8280.605, 8285.697, 8290.61, 8295.341, 8299.883, 8304.234, 8308.398, 8312.374, 8316.165, 8319.774, 8323.211, 8326.4795, 8329.587, 8332.548, 8335.374, 8338.081, 8340.684, 8343.201, 8345.654, 8348.064, 8350.451, 8352.836, 8355.235, 8357.668, 8360.152, 8362.694, 8365.297, 8367.962, 8370.692, 8373.487, 8376.345, 8379.263, 8382.238, 8385.2705, 8388.3545, 8391.488, 8394.669, 8397.892, 8401.151, 8404.441, 8407.758, 8411.095, 8414.447, 8417.809, 8421.175, 8424.541, 8427.907, 8431.27, 8434.626, 8437.979, 8441.329, 8444.68, 8448.034, 8451.394, 8454.761, 8458.139, 8461.53, 8464.9375, 8466.647, 8470.084, 8473.544, 8477.028, 8480.533, 8484.055, 8487.589, 8491.135, 8494.696, 8498.274, 8500.071, 8503.683, 8507.32, 8510.991, 8514.7, 8518.45, 8522.24, 8526.065, 8529.92, 8533.799, 8538.072, 8541.943, 8545.778, 8549.557, 8553.256, 8556.852, 8560.322, 8563.644, 8566.801, 8569.779, 8572.566, 8575.148, 8577.521, 8579.685, 8581.638, 8583.379, 8584.921, 8586.277, 8587.463, 8588.49, 8588.95, 8589.771, 8590.474, 8591.074, 8591.585, 8592.02, 8592.39, 8592.707, 8592.985, 8593.238, 8593.481, 8593.6045, 8593.861, 8594.138, 8594.441, 8594.777, 8595.151, 8595.5625, 8596.011, 8596.493, 8597.009, 8597.554, 8597.836, 8598.417, 8599.017, 8599.629, 8600.246, 8600.859, 8601.46, 8602.043, 8602.607, 8603.153, 8603.681, 8604.19, 8604.692, 8605.192, 8605.698, 8606.222, 8606.776, 8607.382, 8608.052, 8608.803, 8609.642, 8610.578, 8611.622, 8612.779, 8614.051, 8615.439, 8616.946, 8618.569, 8620.303, 8622.139, 8624.072, 8626.093, 8628.189, 8630.352, 8632.567, 8634.825, 8637.118, 8639.4375, 8641.775, 8644.122, 8646.463, 8648.786, 8649.936, 8652.205, 8654.432, 8656.611, 8658.742, 8660.824, 8662.8545, 8664.833, 8666.762, 8668.64, 8669.562, 8671.373, 8673.148, 8674.894, 8676.614, 8678.3125, 8679.989, 8681.647, 8683.287, 8684.909, 8686.514, 8687.309, 8688.887, 8690.445, 8691.9795, 8693.487, 8694.966, 8696.41, 8697.817, 8699.184, 8699.85, 8701.148, 8701.906, 8703.133, 8704.313, 8705.451, 8706.552, 8707.624, 8708.677, 8709.72, 8710.765, 8711.824, 8712.913, 8714.042, 8715.22, 8716.455, 8717.754, 8719.123, 8720.561, 8722.06, 8723.617, 8725.226, 8726.882, 8728.582, 8730.323, 8732.1, 8733.902, 8735.717, 8737.532, 8739.335, 8741.107, 8742.835, 8744.498, 8745.301, 8746.842, 8748.292, 8749.647, 8750.902, 8752.06, 8753.131, 8754.129, 8755.069, 8755.964, 8756.827, 8757.671, 8758.511, 8759.3545, 8760.202, 8761.055, 8761.911, 8762.766, 8763.601, 8764.397, 8765.137, 8765.8, 8766.366, 8766.816, 8767.131, 8767.293, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, -999.0, 8768.357, 8770.835, 8773.3545, 8775.91, 8778.501, 8781.122, 8783.77, 8786.439, 8789.125, 8791.824, 8794.534, 8797.261, 8800.011, 8802.791, 8805.609, 8808.474, 8811.394, 8814.377, 8817.433, 8820.565, 8823.781, 8827.085, 8830.4795, 8833.965, 8837.542, 8841.211, 8844.97, 8848.817, 8852.752, 8856.77, 8860.867, 8865.034, 8869.262, 8873.54, 8877.86, 8882.22, 8886.614, 8891.043, 8895.5, 8899.9795, 8904.476, 8908.98, 8911.234, 8915.74, 8920.236, 8924.716, 8929.17, 8933.595, 8937.989, 8942.351, 8946.676, 8950.966, 8955.22, 8959.438, 8963.622, 8967.77, 8971.88, 8975.951, 8979.982, 8983.97, 8987.906, 8991.787, 8995.605, 8997.491, 9001.218, 9004.886, 9008.499, 9012.061, 9015.581, 9019.069, 9022.535, 9025.987, 9029.424, 9032.845, 9036.249, 9039.636, 9043.005, 9046.3545, 9049.685, 9052.995, 9056.282, 9059.546, 9062.785, 9065.998, 9069.188, 9072.36, 9075.518, 9078.663, 9081.797, 9084.918, 9088.026, 9091.12, 9094.198, 9097.562, 9100.596, 9103.605, 9106.589, 9109.545, 9112.47, 9115.363, 9118.2295, 9121.068, 9123.884, 9126.678, 9129.456, 9132.222, 9134.981, 9137.737, 9140.488, 9143.23, 9145.963, 9148.682, 9151.384, 9154.0625, 9156.716, 9158.03, 9160.64, 9163.224, 9165.785, 9168.327, 9170.854, 9173.368, 9175.874, 9178.376, 9180.879, 9183.392, 9185.919, 9188.471, 9191.051, 9193.665, 9196.32, 9199.021, 9201.773, 9204.583, 9207.456, 9210.398, 9213.416, 9216.514, 9219.697, 9222.974, 9226.341, 9229.797, 9233.339, 9236.961, 9240.662, 9244.438, 9248.286, 9250.236, 9254.184, 9258.189, 9262.245, 9266.341, 9270.47, 9274.622, 9278.791, 9282.966, 9285.054, 9289.225, 9293.383, 9297.522, 9301.636, 9305.718, 9309.768, 9313.78, 9317.754, 9321.6875, 9325.58, 9327.512, 9331.346, 9335.142, 9338.91, 9342.662, 9346.406, 9350.155, 9353.919, 9357.708, 9361.533, 9365.405, 9367.36, 9371.314, 9375.33, 9379.414, 9383.571, 9387.804, 9392.116, 9396.511, 9400.992, 9406.024, 9410.697, 9415.466, 9420.328, 9425.281, 9430.323, 9435.448, 9440.649, 9445.919, 9451.248, 9456.626, 9462.046, 9464.77, 9470.238, 9475.731, 9481.241, 9486.761, 9492.287, 9497.812, 9503.333, 9508.854, 9514.38, 9519.915, 9522.6875, 9528.241, 9533.81, 9539.391, 9544.986, 9550.596, 9556.218, 9561.8545, 9567.504, 9573.167, 9578.847, 9581.692, 9587.3955, 9593.114, 9598.839, 9604.556, 9610.256, 9615.93, 9621.579, 9627.205, 9632.809, 9635.604, 9641.186, 9646.7705, 9652.372, 9658.004, 9663.679, 9669.407, 9675.2, 9681.069, 9687.018, 9693.045, 9699.153, 9705.342, 9711.607, 9717.944, 9724.347, 9730.811, 9737.323, 9743.874, 9750.449, 9757.034, 9760.326, 9766.894, 9773.424, 9779.8955, 9786.291, 9792.598, 9798.803, 9804.8955, 9810.867, 9816.719, 9822.451, 9828.065, 9833.567, 9838.964, 9844.264, 9849.476, 9854.609, 9859.669, 9864.659, 9869.585, 9874.451, 9879.26, 9884.013, 9888.712, 9893.36, 9897.958, 9902.505, 9907.001, 9911.446, 9915.845, 9920.198, 9922.359, 9926.653, 9930.91, 9935.135, 9939.33, 9943.5, 9947.6455, 9951.766, 9955.86, 9959.929, 9961.951, 9965.968, 9969.9375, 9973.851, 9977.697, 9981.471, 9985.164, 9988.772, 9992.289, 9995.713, 9999.37, 10002.597, 10005.7295, 10008.777, 10011.75, 10014.656, 10017.506, 10020.308, 10023.071, 10025.807, 10028.524, 10029.88, 10032.594, 10035.318, 10038.067, 10040.851, 10043.674, 10046.544, 10049.47, 10052.445, 10055.463, 10058.513, 10060.047, 10063.129, 10066.232, 10069.361, 10072.517, 10075.704, 10078.93, 10082.201, 10085.527, 10088.915, 10092.368, 10094.121, 10097.682, 10101.318, 10105.034, 10108.828, 10112.699, 10116.649, 10120.677, 10124.78, 10128.959, 10133.212, 10135.365, 10139.725, 10144.149, 10148.639, 10153.187, 10157.79, 10162.445, 10167.149, 10171.897, 10176.6875, 10181.518, 10183.948, 10188.836, 10193.756, 10198.699, 10203.66, 10208.629, 10213.596, 10218.55, 10223.48, 10228.376, 10233.228, 10238.025, 10242.761, 10247.427, 10252.017, 10256.528, 10260.96, 10265.31, 10269.582, 10273.784, 10277.926, 10282.016, 10286.063, 10290.08, 10294.074, 10298.057, 10302.034, 10306.008, 10309.98, 10313.954, 10317.932, 10319.921, 10323.903, 10327.892, 10331.885, 10335.879, 10339.872, 10343.859, 10347.837, 10351.805, 10356.155, 10360.098, 10364.028, 10367.947, 10371.855, 10375.756, 10379.65, 10383.539, 10387.424, 10391.309, 10395.191, 10397.13, 10401.0, 10404.854, 10408.685, 10412.487, 10416.262, 10420.005, 10423.715, 10427.392, 10431.04, 10434.663, 10438.263, 10441.838, 10445.384, 10448.896, 10452.371, 10455.808, 10459.214, 10462.593, 10465.952, 10469.295, 10470.962, 10474.29, 10477.614, 10480.94, 10484.273, 10487.62, 10490.989, 10494.385, 10497.809, 10501.262, 10502.998, 10506.495, 10510.02, 10513.572, 10517.151, 10520.756, 10524.38, 10528.016, 10531.656, 10535.293, 10538.915, 10542.513, 10544.299, 10547.839, 10551.328, 10554.77, 10558.167, 10561.524, 10564.846, 10568.134, 10571.392, 10574.622, 10577.827, 10581.009, 10584.168, 10587.305, 10590.422, 10593.526, 10596.625, 10599.728, 10602.84, 10605.967, 10607.537, 10610.694, 10613.876, 10617.086, 10620.328, 10623.608, 10626.929, 10630.296, 10633.72, 10637.208, 10640.7705, 10644.409, 10646.257, 10650.01, 10653.839, 10657.739, 10661.701, 10665.712, 10669.757, 10673.824, 10677.91, 10682.009, 10686.116, 10690.228, 10694.337, 10698.435, 10702.515, 10706.568, 10710.598, 10714.601, 10718.58, 10722.537, 10724.901, 10728.825, 10732.732, 10736.626, 10740.5, 10744.347, 10748.158, 10751.927, 10755.6455, 10759.315, 10761.132, 10764.725, 10768.268, 10771.766, 10775.229, 10778.662, 10782.075, 10785.473, 10788.858, 10792.238, 10795.617, 10798.999, 10802.39, 10805.793, 10809.215, 10812.658, 10816.127, 10819.624, 10823.152, 10826.709, 10830.291, 10832.091, 10835.704, 10839.333, 10842.971, 10846.611, 10850.249, 10853.876, 10857.48, 10861.051, 10864.577, 10868.057, 10871.494, 10874.8955, 10878.266, 10881.611, 10884.938, 10888.254, 10891.563, 10894.87, 10898.175, 10901.475, 10904.772, 10908.062, 10911.338, 10914.594, 10917.824, 10921.023, 10924.193, 10927.333, 10930.441, 10933.521, 10936.576, 10939.61, 10941.121, 10944.133, 10947.135, 10950.13, 10953.122}
}
