netcdf file\:/home/walter/TechX/ceres/datasets/WMI_Lear {
  dimensions:
    time = UNLIMITED;   // (180 currently)
  variables:
    double time(time);
      time:units = "seconds since 1970-1-1 0:00:00 0:00";
      time:long_name = "time";
      time:_FillValue = -99999.0;
      time:missing_value = -99999.0;

    float altitude(time);
      altitude:units = "km";
      altitude:long_name = "altitude MSL";
      altitude:_FillValue = -99999.0f;
      altitude:missing_value = -99999.0f;

    float latitude(time);
      latitude:units = "degrees_N";
      latitude:long_name = "latitude";
      latitude:_FillValue = -99999.0f;
      latitude:missing_value = -99999.0f;
      latitude:valid_range = -90.0f, 90.0f;

    float longitude(time);
      longitude:units = "degrees_E";
      longitude:long_name = "longitude";
      longitude:_FillValue = -99999.0f;
      longitude:missing_value = -99999.0f;
      longitude:valid_range = -180.0f, 180.0f;

    float pressure(time);
      pressure:units = "hPa";
      pressure:long_name = "pressure";
      pressure:field_type = "P";
      pressure:_FillValue = -99999.0f;
      pressure:missing_value = -99999.0f;

    float tdry(time);
      tdry:units = "deg_C";
      tdry:long_name = "temperature";
      tdry:field_type = "T";
      tdry:_FillValue = -99999.0f;
      tdry:missing_value = -99999.0f;

    float dp(time);
      dp:units = "deg_C";
      dp:long_name = "dewpoint temperature";
      dp:field_type = "T_d";
      dp:_FillValue = -99999.0f;
      dp:missing_value = -99999.0f;

    float mr(time);
      mr:units = "g/kg";
      mr:long_name = "mixing ratio";
      mr:field_type = "w";
      mr:_FillValue = -99999.0f;
      mr:missing_value = -99999.0f;

    float wspd(time);
      wspd:units = "m/s";
      wspd:long_name = "wind speed";
      wspd:field_type = "wspd";
      wspd:_FillValue = -99999.0f;
      wspd:missing_value = -99999.0f;

    float wdir(time);
      wdir:units = "degrees";
      wdir:long_name = "wind direction";
      wdir:field_type = "wdir";
      wdir:_FillValue = -99999.0f;
      wdir:missing_value = -99999.0f;

    int Drops(time);
      Drops:units = "#";
      Drops:long_name = "Accumulated number of sonde drops";
      Drops:_FillValue = -99999;
      Drops:missing_value = -99999;

  // global attributes:
  :history = "$Id: TrackFile.java,v 1.20 2003/05/07 04:53:23 maclean Exp $";
 data:
time =
  {1.057473013E9, 1.057473019E9, 1.057473029E9, 1.057473039E9, 1.057473049E9, 1.057473059E9, 1.057473069E9, 1.057473079E9, 1.057473089E9, 1.057473099E9, 1.057473109E9, 1.057473119E9, 1.057473129E9, 1.057473139E9, 1.057473149E9, 1.057473159E9, 1.057473169E9, 1.057473179E9, 1.057473189E9, 1.057473199E9, 1.057473209E9, 1.057473219E9, 1.057473229E9, 1.057473239E9, 1.057473249E9, 1.057473259E9, 1.057473269E9, 1.057473279E9, 1.057473289E9, 1.057473299E9, 1.057473309E9, 1.057473319E9, 1.057473329E9, 1.057473339E9, 1.057473349E9, 1.057473359E9, 1.057473369E9, 1.057473379E9, 1.057473389E9, 1.057473399E9, 1.057473409E9, 1.057473419E9, 1.057473429E9, 1.057473439E9, 1.057473449E9, 1.057473459E9, 1.057473469E9, 1.057473479E9, 1.057473489E9, 1.057473499E9, 1.057473509E9, 1.057473519E9, 1.057473529E9, 1.057473539E9, 1.057473549E9, 1.057473559E9, 1.057473569E9, 1.057473579E9, 1.057473589E9, 1.057473599E9, 1.057473609E9, 1.057473619E9, 1.057473629E9, 1.057473639E9, 1.057473649E9, 1.057473659E9, 1.057473669E9, 1.057473679E9, 1.057473689E9, 1.057473699E9, 1.057473709E9, 1.057473719E9, 1.057473729E9, 1.057473739E9, 1.057473749E9, 1.057473759E9, 1.057473769E9, 1.057473779E9, 1.057473789E9, 1.057473799E9, 1.057473809E9, 1.057473819E9, 1.057473829E9, 1.057473839E9, 1.057473849E9, 1.057473859E9, 1.057473869E9, 1.057473879E9, 1.057473889E9, 1.057473899E9, 1.057473909E9, 1.057473919E9, 1.057473929E9, 1.057473939E9, 1.057473949E9, 1.057473959E9, 1.057473969E9, 1.057473979E9, 1.057473989E9, 1.057473999E9, 1.057474009E9, 1.057474019E9, 1.057474029E9, 1.057474039E9, 1.057474049E9, 1.057474059E9, 1.057474069E9, 1.057474079E9, 1.057474089E9, 1.057474099E9, 1.057474109E9, 1.057474119E9, 1.057474129E9, 1.057474139E9, 1.057474149E9, 1.057474159E9, 1.057474169E9, 1.057474179E9, 1.057474189E9, 1.057474199E9, 1.057474209E9, 1.057474219E9, 1.057474229E9, 1.057474239E9, 1.057474249E9, 1.057474259E9, 1.057474269E9, 1.057474279E9, 1.057474289E9, 1.057474299E9, 1.057474309E9, 1.057474319E9, 1.057474329E9, 1.057474339E9, 1.057474349E9, 1.057474359E9, 1.057474369E9, 1.057474379E9, 1.057474389E9, 1.057474399E9, 1.057474409E9, 1.057474419E9, 1.057474429E9, 1.057474439E9, 1.057474449E9, 1.057474459E9, 1.057474469E9, 1.057474479E9, 1.057474489E9, 1.057474499E9, 1.057474509E9, 1.057474519E9, 1.057474529E9, 1.057474539E9, 1.057474549E9, 1.057474559E9, 1.057474569E9, 1.057474579E9, 1.057474589E9, 1.057474599E9, 1.057474609E9, 1.057474619E9, 1.057474629E9, 1.057474639E9, 1.057474649E9, 1.057474659E9, 1.057474669E9, 1.057474679E9, 1.057474689E9, 1.057474699E9, 1.057474709E9, 1.057474719E9, 1.057474729E9, 1.057474739E9, 1.057474749E9, 1.057474759E9, 1.057474769E9, 1.057474779E9, 1.057474789E9, 1.057474799E9}
altitude =
  {0.103, 0.13010001, 0.15210001, 0.18110001, 0.1999, 0.217, 0.228, 0.228, 0.231, 0.2359, 0.2429, 0.25689998, 0.2701, 0.2819, 0.292, 0.3069, 0.3161, 0.3249, 0.331, 0.335, 0.3399, 0.345, 0.349, 0.3511, 0.3539, 0.3569, 0.3591, 0.36089998, 0.3652, 0.3661, 0.37, 0.3719, 0.37489998, 0.37489998, 0.3761, 0.377, 0.378, 0.3801, 0.381, 0.38189998, 0.384, 0.385, 0.3871, 0.38889998, 0.3941, 0.3929, 0.392, 0.392, 0.392, 0.392, 0.4231, 0.5051, 0.612, 0.7251, 0.86990005, 1.0049, 1.1421, 1.2549, 1.471, 1.7291, 1.966, 2.1058998, 2.3158998, 2.485, 2.7011, 2.841, 2.9808998, 3.1018999, 3.191, 3.39, 3.5439, 3.671, 3.778, 3.9621, 4.0709, 4.184, 4.2599, 4.4251003, 4.5839, 4.6939, 4.8881, 5.0271, 5.1401, 5.2388997, 5.4431, 5.5931, 5.729, 5.84, 5.914, 5.979, 6.0981, 6.1692004, 6.2999, 6.4098997, 6.562, 6.68, 6.8409, 6.9561, 7.0229, 7.086, 7.1671, 7.2609, 7.346, 7.4271, 7.5359, 7.6291003, 7.7151003, 7.8291, 7.93, 8.0549, 8.1251, 8.254, 8.357901, 8.5301, 8.6551, 8.847099, 8.918099, 8.92, 8.9261, 8.9559, 9.005, 9.037, 9.1361, 9.2089, 9.315901, 9.3799, 9.5061, 9.586901, 9.6399, 9.6969, 9.746, 9.785, 9.812099, 9.842, 9.9191, 10.002, 10.0721, 10.145, 10.244901, 10.312, 10.3501, 10.3739, 10.378099, 10.3949, 10.465, 10.5379, 10.607, 10.640901, 10.6589, 10.6951, 10.7439, 10.775901, 10.7991, 10.843901, 10.885, 10.935901, 10.977099, 11.0371, 11.0929, 11.135, 11.2051, 11.231, 11.2371, 11.2471, 11.281, 11.3181, 11.3721, 11.401, 11.4541, 11.486099, 11.508, 11.5269, 11.564099, 11.6171, 11.6501, 11.665, 11.679, 11.718, 11.753099, 11.758}
latitude =
  {43.5847, 43.5847, 43.5847, 43.5847, 43.5847, 43.5845, 43.5843, 43.5843, 43.584, 43.5837, 43.5835, 43.5832, 43.583, 43.5832, 43.5833, 43.584, 43.5845, 43.585, 43.5853, 43.5862, 43.5867, 43.5873, 43.5878, 43.5887, 43.5893, 43.59, 43.5908, 43.5913, 43.592, 43.5923, 43.593, 43.5935, 43.5935, 43.5935, 43.5935, 43.5935, 43.5935, 43.5935, 43.5935, 43.5935, 43.5935, 43.5933, 43.5932, 43.5932, 43.5928, 43.5928, 43.5927, 43.5917, 43.5882, 43.5848, 43.5773, 43.5703, 43.5623, 43.5542, 43.5438, 43.5348, 43.5272, 43.5213, 43.513, 43.5065, 43.4997, 43.4948, 43.4865, 43.4798, 43.4707, 43.4633, 43.4543, 43.4445, 43.4373, 43.4235, 43.4118, 43.4022, 43.3947, 43.3808, 43.3698, 43.3573, 43.3493, 43.3353, 43.3235, 43.3153, 43.3, 43.287, 43.2767, 43.2687, 43.2538, 43.243, 43.2322, 43.2207, 43.2113, 43.202, 43.1895, 43.1808, 43.1678, 43.1582, 43.1472, 43.1385, 43.1257, 43.1142, 43.1038, 43.0967, 43.0843, 43.0725, 43.0625, 43.0523, 43.0387, 43.0285, 43.0183, 43.0045, 42.9938, 42.9805, 42.9717, 42.9552, 42.9435, 42.9295, 42.9208, 42.9053, 42.8915, 42.8757, 42.8642, 42.8488, 42.8362, 42.8283, 42.8158, 42.8077, 42.7988, 42.7943, 42.7848, 42.7777, 42.7703, 42.7622, 42.7558, 42.749, 42.7415, 42.7348, 42.7253, 42.7168, 42.7092, 42.7023, 42.6922, 42.683, 42.6752, 42.6682, 42.6573, 42.6488, 42.6373, 42.6283, 42.6182, 42.608, 42.601, 42.5892, 42.5773, 42.5675, 42.5613, 42.549, 42.5363, 42.5268, 42.5177, 42.5065, 42.4962, 42.485, 42.4773, 42.4673, 42.4577, 42.4525, 42.4417, 42.4338, 42.4247, 42.4163, 42.4085, 42.4, 42.3918, 42.384, 42.3738, 42.363, 42.3547, 42.3477, 42.3405, 42.333, 42.326, 42.3207}
longitude =
  {-96.7332, -96.7333, -96.7333, -96.7333, -96.7335, -96.7338, -96.7342, -96.7347, -96.735, -96.7353, -96.7357, -96.7365, -96.737, -96.7373, -96.7375, -96.738, -96.7383, -96.7387, -96.739, -96.7395, -96.7398, -96.7403, -96.7407, -96.7412, -96.7415, -96.742, -96.7425, -96.743, -96.7433, -96.7437, -96.744, -96.7443, -96.7447, -96.7448, -96.745, -96.745, -96.745, -96.745, -96.7448, -96.745, -96.745, -96.7452, -96.7455, -96.7457, -96.7458, -96.7457, -96.7455, -96.745, -96.7427, -96.7405, -96.7358, -96.7318, -96.729, -96.729, -96.7332, -96.7408, -96.7522, -96.7623, -96.7782, -96.7915, -96.8057, -96.8143, -96.8293, -96.8403, -96.8552, -96.8657, -96.8767, -96.8865, -96.893, -96.9047, -96.9143, -96.9223, -96.9285, -96.9402, -96.949, -96.959, -96.9655, -96.9768, -96.986, -96.9923, -97.0037, -97.0137, -97.022, -97.0288, -97.0413, -97.0512, -97.0615, -97.0733, -97.0835, -97.0942, -97.1085, -97.118, -97.1322, -97.1428, -97.1543, -97.1633, -97.1767, -97.1892, -97.2008, -97.2095, -97.2248, -97.2385, -97.2495, -97.2602, -97.2745, -97.2853, -97.296, -97.3102, -97.3203, -97.332, -97.3388, -97.3508, -97.359, -97.3682, -97.3737, -97.3805, -97.3822, -97.3792, -97.374, -97.3625, -97.3482, -97.3365, -97.3117, -97.2913, -97.2688, -97.2567, -97.2302, -97.21, -97.19, -97.168, -97.1495, -97.1288, -97.1085, -97.0927, -97.0683, -97.046, -97.0287, -97.0137, -96.991, -96.9703, -96.9538, -96.939, -96.9167, -96.9, -96.878, -96.8622, -96.845, -96.8277, -96.8155, -96.7942, -96.7727, -96.7548, -96.7443, -96.7233, -96.703, -96.6877, -96.6722, -96.653, -96.6358, -96.617, -96.603, -96.5828, -96.562, -96.5505, -96.5248, -96.5048, -96.4832, -96.4637, -96.4463, -96.4268, -96.4072, -96.3895, -96.3687, -96.3485, -96.3313, -96.3128, -96.2892, -96.2657, -96.2443, -96.2272}
pressure =
  {955.5, 955.5, 955.5, 955.4, 955.5, 955.4, 955.4, 955.5, 955.5, 955.5, 955.4, 955.4, 955.5, 955.4, 955.5, 955.5, 955.5, 955.4, 955.5, 955.5, 955.4, 955.4, 955.4, 955.3, 955.4, 955.3, 955.4, 955.3, 955.3, 955.2, 955.2, 955.3, 955.1, 955.1, 955.1, 955.2, 955.0, 955.1, 955.1, 955.2, 955.0, 955.0, 955.0, 955.0, 955.1, 955.1, 955.0, 954.4, 953.7, 956.5, 949.5, 939.1, 925.9, 912.5, 898.1, 884.0, 869.8, 853.5, 835.6, 808.4, 790.7, 773.9, 757.4, 740.5, 725.9, 713.0, 701.7, 691.7, 679.1, 667.2, 656.1, 644.4, 632.6, 622.9, 614.8, 607.6, 597.8, 586.1, 574.7, 564.0, 554.1, 545.9, 536.8, 526.8, 516.3, 506.7, 498.8, 492.7, 487.9, 482.6, 476.0, 469.7, 463.2, 455.3, 446.3, 438.5, 431.0, 425.6, 421.1, 417.7, 413.8, 408.4, 403.5, 398.9, 393.4, 387.8, 382.9, 378.1, 372.1, 366.7, 361.6, 356.6, 350.3, 342.3, 334.3, 328.3, 326.3, 326.4, 325.8, 323.1, 321.5, 318.3, 315.0, 311.6, 307.3, 302.9, 299.1, 296.1, 294.1, 291.8, 289.7, 288.4, 287.2, 285.2, 282.5, 279.3, 276.2, 272.5, 269.6, 267.8, 265.9, 265.4, 265.0, 264.3, 260.6, 257.8, 256.1, 255.1, 254.0, 252.5, 251.4, 250.1, 249.2, 247.3, 245.7, 244.0, 242.0, 240.4, 238.2, 236.2, 234.8, 234.3, 233.8, 233.3, 232.1, 230.5, 229.0, 227.7, 226.0, 225.1, 224.5, 223.5, 222.3, 220.4, 219.5, 219.0, 217.5, 217.1, 216.6, 215.0}
tdry =
  {21.7, 21.6, 21.6, 21.6, 21.6, 21.6, 21.7, 21.7, 21.6, 21.7, 21.7, 21.6, 21.7, 21.7, 21.7, 21.6, 21.6, 21.6, 21.6, 21.6, 21.6, 21.6, 21.6, 21.6, 21.6, 21.6, 21.6, 21.5, 21.5, 21.5, 21.5, 21.6, 21.8, 22.1, 22.6, 22.7, 22.9, 23.9, 23.8, 23.8, 23.4, 23.1, 22.9, 22.9, 22.8, 22.0, 21.7, 21.6, 21.3, 21.5, 21.9, 22.9, 25.5, 25.4, 25.6, 25.2, 25.3, 26.8, 25.8, 23.0, 21.5, 19.5, 18.3, 16.5, 14.7, 13.0, 11.6, 10.9, 9.6, 8.3, 7.0, 6.3, 6.2, 5.1, 4.2, 5.2, 3.2, 2.5, 0.2, -0.1, -0.9, -1.3, -2.7, -3.8, -4.7, -6.1, -7.2, -7.8, -8.1, -8.2, -8.8, -9.8, -10.1, -10.8, -12.6, -13.9, -15.2, -16.1, -16.7, -16.7, -17.0, -17.4, -18.1, -18.0, -18.6, -19.8, -20.7, -21.9, -22.8, -23.3, -24.1, -23.6, -23.4, -24.3, -25.9, -26.7, -27.0, -26.0, -25.3, -25.0, -25.1, -25.0, -25.6, -25.5, -26.2, -27.4, -28.4, -29.1, -29.5, -30.1, -30.5, -30.7, -30.6, -31.0, -31.6, -32.4, -33.3, -34.1, -35.2, -35.6, -35.6, -35.7, -35.0, -35.3, -35.8, -36.5, -37.0, -37.2, -37.6, -37.7, -38.4, -38.6, -38.9, -39.2, -39.7, -40.3, -41.0, -41.4, -42.1, -42.9, -43.7, -43.7, -43.4, -43.5, -43.8, -43.9, -44.9, -45.4, -45.9, -46.3, -46.2, -46.1, -45.8, -46.2, -46.7, -46.6, -46.3, -47.3, -47.0, -47.8}
dp =
  {14.6, 14.8, 15.0, 15.0, 14.7, 14.8, 14.7, 14.7, 14.7, 14.6, 14.8, 14.8, 14.6, 14.7, 14.9, 14.9, 14.8, 14.8, 14.9, 14.7, 14.5, 14.8, 14.8, 14.6, 14.7, 14.7, 14.7, 14.7, 14.8, 14.8, 14.5, 14.7, 14.7, 15.0, 14.6, 14.8, 14.8, 14.5, 14.5, 15.0, 15.0, 15.3, 15.0, 15.2, 15.2, 15.3, 14.8, 14.7, 14.6, 14.5, 13.5, 12.3, 9.2, 9.2, 7.8, 7.2, 5.9, 4.8, 3.6, 2.6, 2.1, 1.6, 0.8, 0.9, 0.7, 0.5, 0.1, -0.5, -0.8, -1.3, -1.5, -1.2, -2.7, -3.9, -3.8, -6.6, -4.7, -6.2, -7.0, -9.9, -10.0, -7.7, -7.9, -9.0, -10.2, -15.1, -20.9, -25.2, -28.7, -24.7, -15.6, -20.9, -22.6, -26.9, -27.0, -26.4, -26.7, -22.5, -21.4, -19.1, -19.3, -19.1, -20.8, -26.0, -30.2, -33.4, -35.9, -34.7, -33.9, -37.5, -40.4, -42.8, -44.7, -46.1, -47.3, -48.3, -49.1, -48.6, -38.9, -35.9, -39.0, -35.6, -33.9, -34.0, -32.2, -34.0, -32.6, -35.1, -34.7, -33.8, -35.3, -34.4, -33.8, -33.9, -35.1, -36.0, -36.1, -37.1, -37.8, -37.9, -38.4, -38.7, -38.4, -38.4, -39.9, -40.5, -43.0, -43.8, -41.9, -41.8, -42.2, -44.0, -43.6, -42.3, -42.8, -44.5, -44.5, -42.9, -43.9, -45.8, -46.6, -46.8, -46.6, -46.9, -47.2, -47.5, -48.0, -47.7, -47.1, -48.0, -49.2, -50.2, -50.6, -50.8, -50.7, -50.5, -50.9, -51.4, -52.0, -52.4}
mr =
  {11.055769, 11.201944, 11.349853, 11.351062, 11.128641, 11.203137, 11.129827, 11.128641, 11.128641, 11.055769, 11.203137, 11.203137, 11.055769, 11.129827, 11.275681, 11.275681, 11.201944, 11.203137, 11.275681, 11.128641, 10.984494, 11.203137, 11.203137, 11.058125, 11.129827, 11.131013, 11.129827, 11.131013, 11.204332, 11.205525, 10.986835, 11.131013, 11.133385, 11.354693, 11.060481, 11.205525, 11.207915, 10.988006, 10.988006, 11.353482, 11.355904, 11.581177, 11.355904, 11.505643, 11.504416, 11.579942, 11.207915, 11.141697, 11.077006, 10.971639, 10.348013, 9.661859, 7.950433, 8.068699, 7.4484024, 7.2610025, 6.7419267, 6.3607454, 5.968273, 5.745056, 5.6672606, 5.585958, 5.386546, 5.5508513, 5.5815654, 5.6010995, 5.5279236, 5.366694, 5.347529, 5.2460556, 5.2569838, 5.473711, 4.986825, 4.6272783, 4.7243195, 3.8588781, 4.538699, 4.126942, 3.956618, 3.2103732, 3.2421305, 3.9456253, 3.9506748, 3.6925914, 3.4257765, 2.3422258, 1.4507447, 1.000643, 0.7310106, 1.0690732, 2.3920853, 1.5408473, 1.3449391, 0.9265909, 0.93659985, 1.0075681, 0.997171, 1.4771065, 1.6453701, 2.0265286, 2.0107055, 2.07283, 1.8101499, 1.1492449, 0.7867512, 0.58540606, 0.46226594, 0.52794343, 0.5807811, 0.41030017, 0.30788007, 0.2416946, 0.2000159, 0.17526439, 0.15682207, 0.14253215, 0.13082902, 0.13852388, 0.3997753, 0.5478984, 0.40093982, 0.5732165, 0.68617535, 0.68684435, 0.8309723, 0.7065946, 0.82114685, 0.647914, 0.6788977, 0.74815226, 0.64911485, 0.71330476, 0.7601498, 0.75795984, 0.6791397, 0.62754697, 0.62822366, 0.57530516, 0.54129636, 0.53936714, 0.5159421, 0.50111663, 0.5176958, 0.51906806, 0.45034638, 0.42739993, 0.32939526, 0.3031626, 0.37384567, 0.3801111, 0.36576545, 0.30254704, 0.31718123, 0.3678621, 0.35084826, 0.29358077, 0.29600823, 0.35473475, 0.3211587, 0.26266605, 0.24162632, 0.23676056, 0.2426602, 0.23511449, 0.22846782, 0.22237688, 0.21147332, 0.22006279, 0.23730099, 0.21513848, 0.18799192, 0.16815817, 0.16134785, 0.15896918, 0.16150373, 0.1657073, 0.15920949, 0.15038304, 0.14039019, 0.13485637}
wspd =
  {11.7, 11.1, 10.7, 11.2, 10.7, 10.0, 9.8, 10.0, 9.8, 10.9, 9.9, 10.0, 10.0, 9.4, 10.0, 5.7, 3.8, 3.0, 3.0, 2.2, 1.9, 2.8, 1.8, 1.5, 1.1, 1.2, 1.9, 1.4, 2.5, 2.8, 3.3, 7.2, 9.9, 9.8, 10.0, 10.0, 10.0, 10.0, 10.0, 10.0, 10.0, 10.0, 10.0, 10.0, 9.9, 12.6, 14.5, 13.5, 9.8, 8.7, 8.6, 15.4, 22.4, 30.4, 36.1, 34.6, 32.9, 23.1, 16.8, 11.5, 10.7, 11.6, 9.2, 8.6, 9.0, 10.8, 13.8, 14.2, 15.0, 13.3, 13.0, 12.8, 12.4, 15.6, 21.3, 23.0, 25.0, 28.2, 26.4, 24.4, 24.4, 22.3, 21.1, 21.6, 21.5, 18.9, 22.3, 23.1, 24.0, 25.9, 29.6, 29.0, 27.2, 28.0, 26.6, 24.7, 22.4, 19.9, 20.2, 19.3, 20.6, 22.3, 20.7, 20.0, 20.2, 22.2, 22.5, 23.7, 24.2, 23.5, 22.9, 19.7, 17.0, 16.5, 20.2, 28.2, 26.7, 26.5, 27.3, 28.6, 23.8, 25.2, 24.7, 21.2, 19.4, 17.8, 18.6, 16.3, 16.5, 20.0, 20.1, 18.3, 18.4, 19.5, 24.1, 19.5, 18.6, 23.3, 23.8, 24.3, 24.8, 25.5, 22.9, 21.4, 23.3, 22.0, 23.6, 22.4, 24.0, 20.2, 21.0, 17.4, 18.3, 17.6, 20.5, 21.1, 20.7, 16.3, 19.6, 22.8, 23.1, 21.3, 15.5, 13.6, 12.9, 9.1, 10.9, 11.1, 13.9, 16.1, 13.8, 9.0, 10.9, 12.7, 20.5, 23.2, 14.9, 11.1, 13.5, 16.3}
wdir =
  {176.9, 176.9, 176.9, 176.9, 176.9, 195.0, 239.5, 263.0, 241.5, 204.3, 227.5, 241.3, 244.2, 291.1, 331.8, 334.6, 337.3, 338.8, 342.0, 346.7, 347.3, 342.6, 345.6, 353.1, 357.3, 0.2, 346.8, 344.6, 340.1, 341.0, 337.0, 333.1, 320.2, 284.0, 260.8, 259.5, 259.8, 260.0, 260.1, 260.1, 260.1, 255.6, 244.2, 237.4, 214.1, 177.8, 151.6, 151.1, 149.9, 146.4, 133.6, 131.6, 115.8, 99.6, 97.8, 101.7, 103.0, 89.4, 65.5, 43.0, 4.8, 354.3, 7.9, 13.4, 27.1, 9.9, 352.2, 352.4, 356.9, 2.4, 5.4, 6.9, 356.4, 337.6, 330.0, 337.0, 342.4, 340.2, 339.3, 337.5, 333.1, 334.0, 335.8, 332.2, 325.6, 322.5, 316.9, 317.6, 320.7, 324.9, 326.6, 326.2, 328.4, 327.0, 322.0, 314.8, 309.3, 305.6, 307.7, 313.0, 319.2, 322.0, 322.5, 322.2, 321.6, 318.7, 316.6, 315.4, 312.5, 307.4, 303.8, 300.7, 294.4, 278.1, 261.9, 257.4, 247.7, 251.9, 257.9, 260.6, 265.7, 266.7, 266.7, 281.7, 275.9, 264.5, 247.5, 244.9, 239.9, 235.1, 235.9, 240.4, 243.2, 244.7, 236.6, 239.1, 234.0, 222.7, 216.5, 212.7, 212.3, 213.9, 218.6, 224.2, 225.5, 220.3, 214.8, 213.8, 216.1, 216.1, 214.9, 214.1, 214.7, 214.6, 213.8, 213.0, 210.4, 205.2, 204.7, 203.8, 199.5, 197.6, 196.7, 199.9, 203.2, 201.2, 196.6, 192.1, 195.0, 197.1, 196.1, 194.3, 197.2, 195.1, 201.2, 202.6, 202.6, 202.0, 201.2, 202.3}
Drops =
  {0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1}
}
